-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 20 2023 04:45:29

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "ALU_STURCTURE" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of ALU_STURCTURE
entity ALU_STURCTURE is
port (
    S2_S3 : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(7 downto 0);
    F : out std_logic_vector(7 downto 0);
    B : in std_logic_vector(7 downto 0);
    flag_zero : out std_logic;
    A_equal_B : out std_logic;
    B_bigger : out std_logic;
    s2 : in std_logic;
    over_flow : out std_logic;
    carry_out : out std_logic;
    S1 : in std_logic;
    A_bigger : out std_logic;
    CLK : in std_logic);
end ALU_STURCTURE;

-- Architecture of ALU_STURCTURE
-- View name is \INTERFACE\
architecture \INTERFACE\ of ALU_STURCTURE is

signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1884\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1878\ : std_logic;
signal \N__1875\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1818\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1755\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1704\ : std_logic;
signal \N__1701\ : std_logic;
signal \N__1698\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1659\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1650\ : std_logic;
signal \N__1647\ : std_logic;
signal \N__1644\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1614\ : std_logic;
signal \N__1611\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1581\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1566\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1554\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1548\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1539\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1524\ : std_logic;
signal \N__1521\ : std_logic;
signal \N__1518\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1491\ : std_logic;
signal \N__1488\ : std_logic;
signal \N__1485\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1479\ : std_logic;
signal \N__1476\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1452\ : std_logic;
signal \N__1449\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1422\ : std_logic;
signal \N__1419\ : std_logic;
signal \N__1416\ : std_logic;
signal \N__1413\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1392\ : std_logic;
signal \N__1389\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \SYNTHESIZED_WIRE_4_1\ : std_logic;
signal \b2v_inst3.result_reg1_bmZ0Z_0\ : std_logic;
signal \b2v_inst3.result_reg1_amZ0Z_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_3_0_cascade_\ : std_logic;
signal \N_21\ : std_logic;
signal \SYNTHESIZED_WIRE_4_0\ : std_logic;
signal \b2v_inst.A_equal_B_NEZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst.A_equal_B_NEZ0Z_0\ : std_logic;
signal \A_equal_B_c\ : std_logic;
signal \SYNTHESIZED_WIRE_0_4_cascade_\ : std_logic;
signal \b2v_inst4.result_reg2_bmZ0Z_4_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_4\ : std_logic;
signal \SYNTHESIZED_WIRE_0_5_cascade_\ : std_logic;
signal \b2v_inst4.result_reg2_bmZ0Z_5_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_5\ : std_logic;
signal \N_22\ : std_logic;
signal \N_24_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_3\ : std_logic;
signal \b2v_inst4.result_reg2_amZ0Z_4\ : std_logic;
signal \b2v_inst4.result_reg2_amZ0Z_5\ : std_logic;
signal \b2v_inst4.result_reg2_amZ0Z_7_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_7\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \b2v_inst.result_arith_1_1\ : std_logic;
signal \b2v_inst.result_arith_1_cry_0\ : std_logic;
signal \b2v_inst.result_arith_1_cry_1\ : std_logic;
signal \b2v_inst.result_arith_1_3\ : std_logic;
signal \b2v_inst.result_arith_1_cry_2\ : std_logic;
signal b2v_inst_result_arith_1_4 : std_logic;
signal \b2v_inst.result_arith_1_cry_3\ : std_logic;
signal b2v_inst_result_arith_1_5 : std_logic;
signal \b2v_inst.result_arith_1_cry_4\ : std_logic;
signal \b2v_inst.result_arith_1_cry_5\ : std_logic;
signal b2v_inst_result_arith_1_7 : std_logic;
signal \b2v_inst.result_arith_1_cry_6\ : std_logic;
signal \b2v_inst.result_arith_1_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal carry_out_c : std_logic;
signal \b2v_inst.A_c_i_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \b2v_inst.A_c_i_1\ : std_logic;
signal \b2v_inst.B_bigger_cry_0\ : std_logic;
signal \b2v_inst.A_c_i_2\ : std_logic;
signal \b2v_inst.B_bigger_cry_1\ : std_logic;
signal \b2v_inst.A_c_i_3\ : std_logic;
signal \b2v_inst.B_bigger_cry_2\ : std_logic;
signal \b2v_inst.A_c_i_4\ : std_logic;
signal \b2v_inst.B_bigger_cry_3\ : std_logic;
signal \b2v_inst.A_c_i_5\ : std_logic;
signal \b2v_inst.B_bigger_cry_4\ : std_logic;
signal \b2v_inst.A_c_i_6\ : std_logic;
signal \b2v_inst.B_bigger_cry_5\ : std_logic;
signal \b2v_inst.A_c_i_7\ : std_logic;
signal \b2v_inst.B_bigger_cry_6\ : std_logic;
signal \B_bigger_c\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \B_bigger_c_THRU_CO\ : std_logic;
signal \b2v_inst3.result_reg1_amZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst3.result_reg1_bmZ0Z_1\ : std_logic;
signal \SYNTHESIZED_WIRE_3_1\ : std_logic;
signal \b2v_inst3.result_reg1_bmZ0Z_3_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_3_3\ : std_logic;
signal \b2v_inst3.result_reg1_amZ0Z_3\ : std_logic;
signal \b2v_inst.A_equal_B_NEZ0Z_1\ : std_logic;
signal \b2v_inst3.result_reg1_bmZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst3.result_reg1_amZ0Z_2\ : std_logic;
signal \SYNTHESIZED_WIRE_3_2_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_2\ : std_logic;
signal \b2v_inst.A_equal_B_NEZ0Z_3\ : std_logic;
signal \b2v_inst.result_arith_1_2\ : std_logic;
signal \N_23\ : std_logic;
signal s2_c : std_logic;
signal \SYNTHESIZED_WIRE_4_6\ : std_logic;
signal \SYNTHESIZED_WIRE_0_7_cascade_\ : std_logic;
signal \b2v_inst4.result_reg2_bmZ0Z_7\ : std_logic;
signal b2v_inst_result_arith_1_6 : std_logic;
signal \b2v_inst4.result_reg2_amZ0Z_6\ : std_logic;
signal \S2_S3_c_0\ : std_logic;
signal \S2_S3_c_1\ : std_logic;
signal \SYNTHESIZED_WIRE_0_6_cascade_\ : std_logic;
signal \S1_c\ : std_logic;
signal \b2v_inst4.result_reg2_bmZ0Z_6\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_0\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_1\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_2\ : std_logic;
signal \un8_result_arith_cry_3_c_RNIO6R4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_3\ : std_logic;
signal \un8_result_arith_cry_4_c_RNIQ9S4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_4\ : std_logic;
signal \un8_result_arith_cry_5_c_RNISCT4\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_5\ : std_logic;
signal \b2v_inst.un8_result_arith_cry_6\ : std_logic;
signal \un8_result_arith_cry_6_c_RNIK5GH\ : std_logic;
signal \B_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \b2v_inst.B_c_i_0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \A_c_1\ : std_logic;
signal \B_c_1\ : std_logic;
signal \b2v_inst.B_c_i_1\ : std_logic;
signal \b2v_inst.A_bigger_cry_0\ : std_logic;
signal \A_c_2\ : std_logic;
signal \B_c_2\ : std_logic;
signal \b2v_inst.B_c_i_2\ : std_logic;
signal \b2v_inst.A_bigger_cry_1\ : std_logic;
signal \B_c_3\ : std_logic;
signal \A_c_3\ : std_logic;
signal \b2v_inst.B_c_i_3\ : std_logic;
signal \b2v_inst.A_bigger_cry_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \B_c_4\ : std_logic;
signal \b2v_inst.B_c_i_4\ : std_logic;
signal \b2v_inst.A_bigger_cry_3\ : std_logic;
signal \B_c_5\ : std_logic;
signal \A_c_5\ : std_logic;
signal \b2v_inst.B_c_i_5\ : std_logic;
signal \b2v_inst.A_bigger_cry_4\ : std_logic;
signal \B_c_6\ : std_logic;
signal \A_c_6\ : std_logic;
signal \b2v_inst.B_c_i_6\ : std_logic;
signal \b2v_inst.A_bigger_cry_5\ : std_logic;
signal \B_c_7\ : std_logic;
signal \A_c_7\ : std_logic;
signal \b2v_inst.B_c_i_7\ : std_logic;
signal \b2v_inst.A_bigger_cry_6\ : std_logic;
signal \A_bigger_c\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \A_bigger_c_THRU_CO\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(7 downto 0);
signal \B_wire\ : std_logic_vector(7 downto 0);
signal \F_wire\ : std_logic_vector(7 downto 0);
signal \S2_S3_wire\ : std_logic_vector(1 downto 0);
signal carry_out_wire : std_logic;
signal flag_zero_wire : std_logic;
signal \A_equal_B_wire\ : std_logic;
signal \S1_wire\ : std_logic;
signal s2_wire : std_logic;
signal \B_bigger_wire\ : std_logic;
signal over_flow_wire : std_logic;
signal \A_bigger_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \A_wire\ <= A;
    \B_wire\ <= B;
    F <= \F_wire\;
    \S2_S3_wire\ <= S2_S3;
    carry_out <= carry_out_wire;
    flag_zero <= flag_zero_wire;
    A_equal_B <= \A_equal_B_wire\;
    \S1_wire\ <= S1;
    s2_wire <= s2;
    B_bigger <= \B_bigger_wire\;
    over_flow <= over_flow_wire;
    A_bigger <= \A_bigger_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3706\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3708\,
            DIN => \N__3707\,
            DOUT => \N__3706\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3708\,
            PADOUT => \N__3707\,
            PADIN => \N__3706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3697\,
            DIN => \N__3696\,
            DOUT => \N__3695\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3697\,
            PADOUT => \N__3696\,
            PADIN => \N__3695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3688\,
            DIN => \N__3687\,
            DOUT => \N__3686\,
            PACKAGEPIN => \B_wire\(7)
        );

    \B_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3688\,
            PADOUT => \N__3687\,
            PADIN => \N__3686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3679\,
            DIN => \N__3678\,
            DOUT => \N__3677\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3679\,
            PADOUT => \N__3678\,
            PADIN => \N__3677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3670\,
            DIN => \N__3669\,
            DOUT => \N__3668\,
            PACKAGEPIN => \B_wire\(6)
        );

    \B_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3670\,
            PADOUT => \N__3669\,
            PADIN => \N__3668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3661\,
            DIN => \N__3660\,
            DOUT => \N__3659\,
            PACKAGEPIN => \F_wire\(2)
        );

    \F_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3661\,
            PADOUT => \N__3660\,
            PADIN => \N__3659\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1412\
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3652\,
            DIN => \N__3651\,
            DOUT => \N__3650\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3652\,
            PADOUT => \N__3651\,
            PADIN => \N__3650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3643\,
            DIN => \N__3642\,
            DOUT => \N__3641\,
            PACKAGEPIN => \B_wire\(2)
        );

    \B_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3643\,
            PADOUT => \N__3642\,
            PADIN => \N__3641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3634\,
            DIN => \N__3633\,
            DOUT => \N__3632\,
            PACKAGEPIN => \F_wire\(5)
        );

    \F_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3634\,
            PADOUT => \N__3633\,
            PADIN => \N__3632\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1409\
        );

    \S2_S3_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3625\,
            DIN => \N__3624\,
            DOUT => \N__3623\,
            PACKAGEPIN => \S2_S3_wire\(0)
        );

    \S2_S3_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3625\,
            PADOUT => \N__3624\,
            PADIN => \N__3623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \S2_S3_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \carry_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3616\,
            DIN => \N__3615\,
            DOUT => \N__3614\,
            PACKAGEPIN => carry_out_wire
        );

    \carry_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3616\,
            PADOUT => \N__3615\,
            PADIN => \N__3614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \flag_zero_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3607\,
            DIN => \N__3606\,
            DOUT => \N__3605\,
            PACKAGEPIN => flag_zero_wire
        );

    \flag_zero_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3607\,
            PADOUT => \N__3606\,
            PADIN => \N__3605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1392\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3598\,
            DIN => \N__3597\,
            DOUT => \N__3596\,
            PACKAGEPIN => \F_wire\(1)
        );

    \F_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3598\,
            PADOUT => \N__3597\,
            PADIN => \N__3596\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1413\
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3589\,
            DIN => \N__3588\,
            DOUT => \N__3587\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3589\,
            PADOUT => \N__3588\,
            PADIN => \N__3587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3580\,
            DIN => \N__3579\,
            DOUT => \N__3578\,
            PACKAGEPIN => \B_wire\(5)
        );

    \B_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3580\,
            PADOUT => \N__3579\,
            PADIN => \N__3578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3571\,
            DIN => \N__3570\,
            DOUT => \N__3569\,
            PACKAGEPIN => \F_wire\(4)
        );

    \F_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3571\,
            PADOUT => \N__3570\,
            PADIN => \N__3569\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1411\
        );

    \A_equal_B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3562\,
            DIN => \N__3561\,
            DOUT => \N__3560\,
            PACKAGEPIN => \A_equal_B_wire\
        );

    \A_equal_B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3562\,
            PADOUT => \N__3561\,
            PADIN => \N__3560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \S1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3553\,
            DIN => \N__3552\,
            DOUT => \N__3551\,
            PACKAGEPIN => \S1_wire\
        );

    \S1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3553\,
            PADOUT => \N__3552\,
            PADIN => \N__3551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \S1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3544\,
            DIN => \N__3543\,
            DOUT => \N__3542\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3544\,
            PADOUT => \N__3543\,
            PADIN => \N__3542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3535\,
            DIN => \N__3534\,
            DOUT => \N__3533\,
            PACKAGEPIN => \B_wire\(1)
        );

    \B_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3535\,
            PADOUT => \N__3534\,
            PADIN => \N__3533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3526\,
            DIN => \N__3525\,
            DOUT => \N__3524\,
            PACKAGEPIN => \F_wire\(0)
        );

    \F_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3526\,
            PADOUT => \N__3525\,
            PADIN => \N__3524\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1411\
        );

    \s2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3517\,
            DIN => \N__3516\,
            DOUT => \N__3515\,
            PACKAGEPIN => s2_wire
        );

    \s2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3517\,
            PADOUT => \N__3516\,
            PADIN => \N__3515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => s2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_bigger_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3508\,
            DIN => \N__3507\,
            DOUT => \N__3506\,
            PACKAGEPIN => \B_bigger_wire\
        );

    \B_bigger_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3508\,
            PADOUT => \N__3507\,
            PADIN => \N__3506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1731\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3499\,
            DIN => \N__3498\,
            DOUT => \N__3497\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3499\,
            PADOUT => \N__3498\,
            PADIN => \N__3497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3490\,
            DIN => \N__3489\,
            DOUT => \N__3488\,
            PACKAGEPIN => \B_wire\(4)
        );

    \B_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3490\,
            PADOUT => \N__3489\,
            PADIN => \N__3488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \over_flow_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3481\,
            DIN => \N__3480\,
            DOUT => \N__3479\,
            PACKAGEPIN => over_flow_wire
        );

    \over_flow_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3481\,
            PADOUT => \N__3480\,
            PADIN => \N__3479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3472\,
            DIN => \N__3471\,
            DOUT => \N__3470\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3472\,
            PADOUT => \N__3471\,
            PADIN => \N__3470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3463\,
            DIN => \N__3462\,
            DOUT => \N__3461\,
            PACKAGEPIN => \B_wire\(0)
        );

    \B_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3463\,
            PADOUT => \N__3462\,
            PADIN => \N__3461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3454\,
            DIN => \N__3453\,
            DOUT => \N__3452\,
            PACKAGEPIN => \F_wire\(7)
        );

    \F_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3454\,
            PADOUT => \N__3453\,
            PADIN => \N__3452\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1605\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1410\
        );

    \A_bigger_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3445\,
            DIN => \N__3444\,
            DOUT => \N__3443\,
            PACKAGEPIN => \A_bigger_wire\
        );

    \A_bigger_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3445\,
            PADOUT => \N__3444\,
            PADIN => \N__3443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3436\,
            DIN => \N__3435\,
            DOUT => \N__3434\,
            PACKAGEPIN => \F_wire\(3)
        );

    \F_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3436\,
            PADOUT => \N__3435\,
            PADIN => \N__3434\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1509\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1412\
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3427\,
            DIN => \N__3426\,
            DOUT => \N__3425\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3427\,
            PADOUT => \N__3426\,
            PADIN => \N__3425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3418\,
            DIN => \N__3417\,
            DOUT => \N__3416\,
            PACKAGEPIN => \B_wire\(3)
        );

    \B_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3418\,
            PADOUT => \N__3417\,
            PADIN => \N__3416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3409\,
            DIN => \N__3408\,
            DOUT => \N__3407\,
            PACKAGEPIN => \F_wire\(6)
        );

    \F_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__3409\,
            PADOUT => \N__3408\,
            PADIN => \N__3407\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1755\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1410\
        );

    \S2_S3_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3400\,
            DIN => \N__3399\,
            DOUT => \N__3398\,
            PACKAGEPIN => \S2_S3_wire\(1)
        );

    \S2_S3_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3400\,
            PADOUT => \N__3399\,
            PADIN => \N__3398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \S2_S3_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__786\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3370\
        );

    \I__785\ : InMux
    port map (
            O => \N__3380\,
            I => \N__3370\
        );

    \I__784\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3370\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__3378\,
            I => \N__3366\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \N__3363\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3370\,
            I => \N__3360\
        );

    \I__780\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3357\
        );

    \I__779\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3354\
        );

    \I__778\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3351\
        );

    \I__777\ : Span4Mux_s1_h
    port map (
            O => \N__3360\,
            I => \N__3344\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3357\,
            I => \N__3344\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3354\,
            I => \N__3344\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3351\,
            I => \N__3341\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__3344\,
            I => \N__3337\
        );

    \I__772\ : Span4Mux_v
    port map (
            O => \N__3341\,
            I => \N__3334\
        );

    \I__771\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3331\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__3337\,
            I => \A_c_4\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3334\,
            I => \A_c_4\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3331\,
            I => \A_c_4\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__3324\,
            I => \N__3319\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__3323\,
            I => \N__3316\
        );

    \I__765\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3311\
        );

    \I__764\ : InMux
    port map (
            O => \N__3319\,
            I => \N__3311\
        );

    \I__763\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3308\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3311\,
            I => \N__3303\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3308\,
            I => \N__3300\
        );

    \I__760\ : InMux
    port map (
            O => \N__3307\,
            I => \N__3297\
        );

    \I__759\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3294\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__3303\,
            I => \N__3289\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__3300\,
            I => \N__3289\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__3297\,
            I => \N__3286\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3294\,
            I => \B_c_4\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__3289\,
            I => \B_c_4\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__3286\,
            I => \B_c_4\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__751\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3272\
        );

    \I__750\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3269\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3272\,
            I => \b2v_inst.B_c_i_4\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3269\,
            I => \b2v_inst.B_c_i_4\
        );

    \I__747\ : InMux
    port map (
            O => \N__3264\,
            I => \N__3258\
        );

    \I__746\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3258\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3258\,
            I => \N__3253\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__3257\,
            I => \N__3249\
        );

    \I__743\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3246\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__3253\,
            I => \N__3243\
        );

    \I__741\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3240\
        );

    \I__740\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3237\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3246\,
            I => \N__3234\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__3243\,
            I => \B_c_5\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3240\,
            I => \B_c_5\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3237\,
            I => \B_c_5\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__3234\,
            I => \B_c_5\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__3225\,
            I => \N__3218\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3224\,
            I => \N__3214\
        );

    \I__732\ : InMux
    port map (
            O => \N__3223\,
            I => \N__3211\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__3222\,
            I => \N__3208\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__3221\,
            I => \N__3205\
        );

    \I__729\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3200\
        );

    \I__728\ : InMux
    port map (
            O => \N__3217\,
            I => \N__3200\
        );

    \I__727\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3196\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3211\,
            I => \N__3193\
        );

    \I__725\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3190\
        );

    \I__724\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3187\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3200\,
            I => \N__3184\
        );

    \I__722\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3181\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3196\,
            I => \N__3178\
        );

    \I__720\ : Span4Mux_s3_h
    port map (
            O => \N__3193\,
            I => \N__3175\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3190\,
            I => \N__3170\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3187\,
            I => \N__3170\
        );

    \I__717\ : Span4Mux_s3_h
    port map (
            O => \N__3184\,
            I => \N__3167\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3181\,
            I => \N__3164\
        );

    \I__715\ : Span4Mux_s3_h
    port map (
            O => \N__3178\,
            I => \N__3161\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__3175\,
            I => \N__3158\
        );

    \I__713\ : Span12Mux_s3_h
    port map (
            O => \N__3170\,
            I => \N__3155\
        );

    \I__712\ : Span4Mux_v
    port map (
            O => \N__3167\,
            I => \N__3150\
        );

    \I__711\ : Span4Mux_s3_h
    port map (
            O => \N__3164\,
            I => \N__3150\
        );

    \I__710\ : Span4Mux_v
    port map (
            O => \N__3161\,
            I => \N__3147\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__3158\,
            I => \A_c_5\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__3155\,
            I => \A_c_5\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3150\,
            I => \A_c_5\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3147\,
            I => \A_c_5\
        );

    \I__705\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3134\
        );

    \I__704\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3131\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3134\,
            I => \b2v_inst.B_c_i_5\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3131\,
            I => \b2v_inst.B_c_i_5\
        );

    \I__701\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3118\
        );

    \I__700\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3118\
        );

    \I__699\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3115\
        );

    \I__698\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3112\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3118\,
            I => \N__3104\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3115\,
            I => \N__3104\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3112\,
            I => \N__3104\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3111\,
            I => \N__3101\
        );

    \I__693\ : Span4Mux_v
    port map (
            O => \N__3104\,
            I => \N__3098\
        );

    \I__692\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3095\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__3098\,
            I => \B_c_6\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3095\,
            I => \B_c_6\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__3090\,
            I => \N__3085\
        );

    \I__688\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3075\
        );

    \I__687\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3075\
        );

    \I__686\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3075\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__3084\,
            I => \N__3072\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3083\,
            I => \N__3069\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \N__3066\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3075\,
            I => \N__3063\
        );

    \I__681\ : InMux
    port map (
            O => \N__3072\,
            I => \N__3060\
        );

    \I__680\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3057\
        );

    \I__679\ : InMux
    port map (
            O => \N__3066\,
            I => \N__3054\
        );

    \I__678\ : Span4Mux_h
    port map (
            O => \N__3063\,
            I => \N__3047\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3060\,
            I => \N__3047\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3057\,
            I => \N__3047\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3054\,
            I => \N__3044\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__3047\,
            I => \N__3040\
        );

    \I__673\ : Span4Mux_v
    port map (
            O => \N__3044\,
            I => \N__3037\
        );

    \I__672\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3034\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__3040\,
            I => \A_c_6\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__3037\,
            I => \A_c_6\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3034\,
            I => \A_c_6\
        );

    \I__668\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3023\
        );

    \I__667\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3020\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3023\,
            I => \b2v_inst.B_c_i_6\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3020\,
            I => \b2v_inst.B_c_i_6\
        );

    \I__664\ : InMux
    port map (
            O => \N__3015\,
            I => \N__3007\
        );

    \I__663\ : InMux
    port map (
            O => \N__3014\,
            I => \N__3007\
        );

    \I__662\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3004\
        );

    \I__661\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3001\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3007\,
            I => \N__2997\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3004\,
            I => \N__2994\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3001\,
            I => \N__2991\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__3000\,
            I => \N__2987\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__2997\,
            I => \N__2984\
        );

    \I__655\ : Span4Mux_h
    port map (
            O => \N__2994\,
            I => \N__2981\
        );

    \I__654\ : Span4Mux_h
    port map (
            O => \N__2991\,
            I => \N__2978\
        );

    \I__653\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2975\
        );

    \I__652\ : InMux
    port map (
            O => \N__2987\,
            I => \N__2972\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__2984\,
            I => \N__2969\
        );

    \I__650\ : Span4Mux_v
    port map (
            O => \N__2981\,
            I => \N__2966\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__2978\,
            I => \N__2959\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__2975\,
            I => \N__2959\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2959\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__2969\,
            I => \B_c_7\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__2966\,
            I => \B_c_7\
        );

    \I__644\ : Odrv12
    port map (
            O => \N__2959\,
            I => \B_c_7\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__642\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2941\
        );

    \I__641\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2941\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__2947\,
            I => \N__2938\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__2946\,
            I => \N__2934\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2931\
        );

    \I__637\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2928\
        );

    \I__636\ : InMux
    port map (
            O => \N__2937\,
            I => \N__2925\
        );

    \I__635\ : InMux
    port map (
            O => \N__2934\,
            I => \N__2922\
        );

    \I__634\ : Span4Mux_h
    port map (
            O => \N__2931\,
            I => \N__2917\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__2928\,
            I => \N__2917\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__2925\,
            I => \N__2914\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__2922\,
            I => \N__2911\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__2917\,
            I => \N__2907\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__2914\,
            I => \N__2902\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__2911\,
            I => \N__2902\
        );

    \I__627\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2899\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__2907\,
            I => \A_c_7\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__2902\,
            I => \A_c_7\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__2899\,
            I => \A_c_7\
        );

    \I__623\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__2889\,
            I => \b2v_inst.B_c_i_7\
        );

    \I__621\ : InMux
    port map (
            O => \N__2886\,
            I => \bfn_2_13_0_\
        );

    \I__620\ : IoInMux
    port map (
            O => \N__2883\,
            I => \N__2880\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__618\ : Span4Mux_s3_v
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__2874\,
            I => \A_bigger_c_THRU_CO\
        );

    \I__616\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__2868\,
            I => \un8_result_arith_cry_4_c_RNIQ9S4\
        );

    \I__614\ : InMux
    port map (
            O => \N__2865\,
            I => \b2v_inst.un8_result_arith_cry_4\
        );

    \I__613\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2859\,
            I => \un8_result_arith_cry_5_c_RNISCT4\
        );

    \I__611\ : InMux
    port map (
            O => \N__2856\,
            I => \b2v_inst.un8_result_arith_cry_5\
        );

    \I__610\ : InMux
    port map (
            O => \N__2853\,
            I => \b2v_inst.un8_result_arith_cry_6\
        );

    \I__609\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__2847\,
            I => \un8_result_arith_cry_6_c_RNIK5GH\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__2844\,
            I => \N__2839\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__2843\,
            I => \N__2835\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__2842\,
            I => \N__2832\
        );

    \I__604\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2828\
        );

    \I__603\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2823\
        );

    \I__602\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2823\
        );

    \I__601\ : InMux
    port map (
            O => \N__2832\,
            I => \N__2820\
        );

    \I__600\ : InMux
    port map (
            O => \N__2831\,
            I => \N__2817\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__2828\,
            I => \N__2814\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__2823\,
            I => \N__2811\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__2820\,
            I => \N__2806\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__2817\,
            I => \N__2806\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__2814\,
            I => \N__2798\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__2811\,
            I => \N__2798\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__2806\,
            I => \N__2798\
        );

    \I__592\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2795\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__2798\,
            I => \B_c_0\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__2795\,
            I => \B_c_0\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__588\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2775\
        );

    \I__587\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2775\
        );

    \I__586\ : InMux
    port map (
            O => \N__2785\,
            I => \N__2775\
        );

    \I__585\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2772\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__2783\,
            I => \N__2767\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__2782\,
            I => \N__2764\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2775\,
            I => \N__2761\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__2772\,
            I => \N__2758\
        );

    \I__580\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2755\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__2770\,
            I => \N__2752\
        );

    \I__578\ : InMux
    port map (
            O => \N__2767\,
            I => \N__2748\
        );

    \I__577\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2745\
        );

    \I__576\ : Span4Mux_s2_h
    port map (
            O => \N__2761\,
            I => \N__2741\
        );

    \I__575\ : Span4Mux_s2_h
    port map (
            O => \N__2758\,
            I => \N__2738\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2755\,
            I => \N__2735\
        );

    \I__573\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2732\
        );

    \I__572\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2729\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__2748\,
            I => \N__2726\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__2745\,
            I => \N__2723\
        );

    \I__569\ : InMux
    port map (
            O => \N__2744\,
            I => \N__2720\
        );

    \I__568\ : Span4Mux_v
    port map (
            O => \N__2741\,
            I => \N__2715\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__2738\,
            I => \N__2715\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__2735\,
            I => \N__2710\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2732\,
            I => \N__2710\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__2729\,
            I => \N__2707\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__2726\,
            I => \N__2700\
        );

    \I__562\ : Span4Mux_s2_h
    port map (
            O => \N__2723\,
            I => \N__2700\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2700\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__2715\,
            I => \N__2697\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__2710\,
            I => \N__2692\
        );

    \I__558\ : Span4Mux_s2_h
    port map (
            O => \N__2707\,
            I => \N__2692\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__2700\,
            I => \N__2689\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__2697\,
            I => \A_c_0\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__2692\,
            I => \A_c_0\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__2689\,
            I => \A_c_0\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__2682\,
            I => \N__2678\
        );

    \I__552\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2675\
        );

    \I__551\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2672\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2675\,
            I => \b2v_inst.B_c_i_0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2672\,
            I => \b2v_inst.B_c_i_0\
        );

    \I__548\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2658\
        );

    \I__547\ : InMux
    port map (
            O => \N__2666\,
            I => \N__2658\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__2665\,
            I => \N__2654\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__2664\,
            I => \N__2651\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__2663\,
            I => \N__2647\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2658\,
            I => \N__2644\
        );

    \I__542\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2640\
        );

    \I__541\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2637\
        );

    \I__540\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2634\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__2650\,
            I => \N__2631\
        );

    \I__538\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2628\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__2644\,
            I => \N__2625\
        );

    \I__536\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2622\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__2640\,
            I => \N__2617\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2637\,
            I => \N__2617\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2634\,
            I => \N__2614\
        );

    \I__532\ : InMux
    port map (
            O => \N__2631\,
            I => \N__2611\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__2628\,
            I => \N__2608\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__2625\,
            I => \N__2605\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__2622\,
            I => \N__2602\
        );

    \I__528\ : Span4Mux_v
    port map (
            O => \N__2617\,
            I => \N__2595\
        );

    \I__527\ : Span4Mux_s2_h
    port map (
            O => \N__2614\,
            I => \N__2595\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__2611\,
            I => \N__2595\
        );

    \I__525\ : Span4Mux_v
    port map (
            O => \N__2608\,
            I => \N__2592\
        );

    \I__524\ : IoSpan4Mux
    port map (
            O => \N__2605\,
            I => \N__2587\
        );

    \I__523\ : IoSpan4Mux
    port map (
            O => \N__2602\,
            I => \N__2587\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__2595\,
            I => \N__2584\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__2592\,
            I => \A_c_1\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__2587\,
            I => \A_c_1\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__2584\,
            I => \A_c_1\
        );

    \I__518\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2571\
        );

    \I__517\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2568\
        );

    \I__516\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2565\
        );

    \I__515\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2562\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2571\,
            I => \N__2559\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2568\,
            I => \N__2556\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2565\,
            I => \N__2553\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2562\,
            I => \N__2550\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__2559\,
            I => \N__2544\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__2556\,
            I => \N__2544\
        );

    \I__508\ : Span4Mux_v
    port map (
            O => \N__2553\,
            I => \N__2539\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__2550\,
            I => \N__2539\
        );

    \I__506\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2536\
        );

    \I__505\ : Odrv4
    port map (
            O => \N__2544\,
            I => \B_c_1\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__2539\,
            I => \B_c_1\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2536\,
            I => \B_c_1\
        );

    \I__502\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2525\
        );

    \I__501\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2522\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2525\,
            I => \b2v_inst.B_c_i_1\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2522\,
            I => \b2v_inst.B_c_i_1\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__2517\,
            I => \N__2512\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__2516\,
            I => \N__2508\
        );

    \I__496\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2505\
        );

    \I__495\ : InMux
    port map (
            O => \N__2512\,
            I => \N__2502\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__2511\,
            I => \N__2498\
        );

    \I__493\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2495\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2505\,
            I => \N__2489\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2502\,
            I => \N__2486\
        );

    \I__490\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2483\
        );

    \I__489\ : InMux
    port map (
            O => \N__2498\,
            I => \N__2480\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2495\,
            I => \N__2477\
        );

    \I__487\ : InMux
    port map (
            O => \N__2494\,
            I => \N__2470\
        );

    \I__486\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2470\
        );

    \I__485\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2470\
        );

    \I__484\ : Span4Mux_s1_h
    port map (
            O => \N__2489\,
            I => \N__2461\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__2486\,
            I => \N__2461\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2483\,
            I => \N__2461\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2480\,
            I => \N__2461\
        );

    \I__480\ : Sp12to4
    port map (
            O => \N__2477\,
            I => \N__2456\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2470\,
            I => \N__2456\
        );

    \I__478\ : Span4Mux_v
    port map (
            O => \N__2461\,
            I => \N__2453\
        );

    \I__477\ : Odrv12
    port map (
            O => \N__2456\,
            I => \A_c_2\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__2453\,
            I => \A_c_2\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__2448\,
            I => \N__2443\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__2447\,
            I => \N__2440\
        );

    \I__473\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2437\
        );

    \I__472\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2431\
        );

    \I__471\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2431\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2437\,
            I => \N__2428\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__2436\,
            I => \N__2425\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2431\,
            I => \N__2422\
        );

    \I__467\ : Span4Mux_h
    port map (
            O => \N__2428\,
            I => \N__2418\
        );

    \I__466\ : InMux
    port map (
            O => \N__2425\,
            I => \N__2415\
        );

    \I__465\ : Span4Mux_h
    port map (
            O => \N__2422\,
            I => \N__2412\
        );

    \I__464\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2409\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__2418\,
            I => \N__2406\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2415\,
            I => \N__2403\
        );

    \I__461\ : Sp12to4
    port map (
            O => \N__2412\,
            I => \N__2398\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2409\,
            I => \N__2398\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__2406\,
            I => \B_c_2\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__2403\,
            I => \B_c_2\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__2398\,
            I => \B_c_2\
        );

    \I__456\ : InMux
    port map (
            O => \N__2391\,
            I => \N__2387\
        );

    \I__455\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2384\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2387\,
            I => \b2v_inst.B_c_i_2\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2384\,
            I => \b2v_inst.B_c_i_2\
        );

    \I__452\ : InMux
    port map (
            O => \N__2379\,
            I => \N__2374\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__2378\,
            I => \N__2371\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__2377\,
            I => \N__2368\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2374\,
            I => \N__2364\
        );

    \I__448\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2361\
        );

    \I__447\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2355\
        );

    \I__446\ : InMux
    port map (
            O => \N__2367\,
            I => \N__2355\
        );

    \I__445\ : Span4Mux_v
    port map (
            O => \N__2364\,
            I => \N__2350\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2361\,
            I => \N__2350\
        );

    \I__443\ : InMux
    port map (
            O => \N__2360\,
            I => \N__2347\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2355\,
            I => \N__2344\
        );

    \I__441\ : Span4Mux_v
    port map (
            O => \N__2350\,
            I => \N__2341\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2347\,
            I => \N__2338\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__2344\,
            I => \B_c_3\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__2341\,
            I => \B_c_3\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__2338\,
            I => \B_c_3\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__2331\,
            I => \N__2325\
        );

    \I__435\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2315\
        );

    \I__434\ : InMux
    port map (
            O => \N__2329\,
            I => \N__2315\
        );

    \I__433\ : InMux
    port map (
            O => \N__2328\,
            I => \N__2315\
        );

    \I__432\ : InMux
    port map (
            O => \N__2325\,
            I => \N__2312\
        );

    \I__431\ : InMux
    port map (
            O => \N__2324\,
            I => \N__2308\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__2323\,
            I => \N__2305\
        );

    \I__429\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2302\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2315\,
            I => \N__2297\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2312\,
            I => \N__2297\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__2311\,
            I => \N__2294\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2308\,
            I => \N__2291\
        );

    \I__424\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2288\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2302\,
            I => \N__2284\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__2297\,
            I => \N__2281\
        );

    \I__421\ : InMux
    port map (
            O => \N__2294\,
            I => \N__2278\
        );

    \I__420\ : Span4Mux_s2_h
    port map (
            O => \N__2291\,
            I => \N__2273\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2288\,
            I => \N__2273\
        );

    \I__418\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2270\
        );

    \I__417\ : Span4Mux_s3_h
    port map (
            O => \N__2284\,
            I => \N__2267\
        );

    \I__416\ : IoSpan4Mux
    port map (
            O => \N__2281\,
            I => \N__2262\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2278\,
            I => \N__2262\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__2273\,
            I => \N__2259\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2270\,
            I => \N__2256\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__2267\,
            I => \N__2251\
        );

    \I__411\ : Span4Mux_s3_h
    port map (
            O => \N__2262\,
            I => \N__2251\
        );

    \I__410\ : IoSpan4Mux
    port map (
            O => \N__2259\,
            I => \N__2248\
        );

    \I__409\ : Span4Mux_s3_h
    port map (
            O => \N__2256\,
            I => \N__2245\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__2251\,
            I => \N__2242\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__2248\,
            I => \A_c_3\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__2245\,
            I => \A_c_3\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__2242\,
            I => \A_c_3\
        );

    \I__404\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2231\
        );

    \I__403\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2228\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2231\,
            I => \b2v_inst.B_c_i_3\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2228\,
            I => \b2v_inst.B_c_i_3\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__2223\,
            I => \SYNTHESIZED_WIRE_0_7_cascade_\
        );

    \I__399\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2217\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2217\,
            I => \b2v_inst4.result_reg2_bmZ0Z_7\
        );

    \I__397\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2211\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2211\,
            I => b2v_inst_result_arith_1_6
        );

    \I__395\ : InMux
    port map (
            O => \N__2208\,
            I => \N__2205\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2205\,
            I => \b2v_inst4.result_reg2_amZ0Z_6\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__2202\,
            I => \N__2198\
        );

    \I__392\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2180\
        );

    \I__391\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2180\
        );

    \I__390\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2175\
        );

    \I__389\ : InMux
    port map (
            O => \N__2196\,
            I => \N__2175\
        );

    \I__388\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2166\
        );

    \I__387\ : InMux
    port map (
            O => \N__2194\,
            I => \N__2166\
        );

    \I__386\ : InMux
    port map (
            O => \N__2193\,
            I => \N__2166\
        );

    \I__385\ : InMux
    port map (
            O => \N__2192\,
            I => \N__2166\
        );

    \I__384\ : InMux
    port map (
            O => \N__2191\,
            I => \N__2163\
        );

    \I__383\ : InMux
    port map (
            O => \N__2190\,
            I => \N__2152\
        );

    \I__382\ : InMux
    port map (
            O => \N__2189\,
            I => \N__2152\
        );

    \I__381\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2152\
        );

    \I__380\ : InMux
    port map (
            O => \N__2187\,
            I => \N__2152\
        );

    \I__379\ : InMux
    port map (
            O => \N__2186\,
            I => \N__2152\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2185\,
            I => \N__2147\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2180\,
            I => \N__2139\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2175\,
            I => \N__2139\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2166\,
            I => \N__2139\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2163\,
            I => \N__2134\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2152\,
            I => \N__2134\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2151\,
            I => \N__2130\
        );

    \I__371\ : InMux
    port map (
            O => \N__2150\,
            I => \N__2125\
        );

    \I__370\ : InMux
    port map (
            O => \N__2147\,
            I => \N__2125\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__2146\,
            I => \N__2122\
        );

    \I__368\ : Span4Mux_v
    port map (
            O => \N__2139\,
            I => \N__2117\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__2134\,
            I => \N__2114\
        );

    \I__366\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2109\
        );

    \I__365\ : InMux
    port map (
            O => \N__2130\,
            I => \N__2109\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2125\,
            I => \N__2106\
        );

    \I__363\ : InMux
    port map (
            O => \N__2122\,
            I => \N__2103\
        );

    \I__362\ : InMux
    port map (
            O => \N__2121\,
            I => \N__2098\
        );

    \I__361\ : InMux
    port map (
            O => \N__2120\,
            I => \N__2098\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__2117\,
            I => \S2_S3_c_0\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__2114\,
            I => \S2_S3_c_0\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2109\,
            I => \S2_S3_c_0\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__2106\,
            I => \S2_S3_c_0\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2103\,
            I => \S2_S3_c_0\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2098\,
            I => \S2_S3_c_0\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2085\,
            I => \N__2075\
        );

    \I__353\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2065\
        );

    \I__352\ : InMux
    port map (
            O => \N__2083\,
            I => \N__2060\
        );

    \I__351\ : InMux
    port map (
            O => \N__2082\,
            I => \N__2060\
        );

    \I__350\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2055\
        );

    \I__349\ : InMux
    port map (
            O => \N__2080\,
            I => \N__2055\
        );

    \I__348\ : InMux
    port map (
            O => \N__2079\,
            I => \N__2044\
        );

    \I__347\ : InMux
    port map (
            O => \N__2078\,
            I => \N__2044\
        );

    \I__346\ : InMux
    port map (
            O => \N__2075\,
            I => \N__2044\
        );

    \I__345\ : InMux
    port map (
            O => \N__2074\,
            I => \N__2044\
        );

    \I__344\ : InMux
    port map (
            O => \N__2073\,
            I => \N__2044\
        );

    \I__343\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2033\
        );

    \I__342\ : InMux
    port map (
            O => \N__2071\,
            I => \N__2033\
        );

    \I__341\ : InMux
    port map (
            O => \N__2070\,
            I => \N__2033\
        );

    \I__340\ : InMux
    port map (
            O => \N__2069\,
            I => \N__2033\
        );

    \I__339\ : InMux
    port map (
            O => \N__2068\,
            I => \N__2033\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2065\,
            I => \N__2024\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2060\,
            I => \N__2024\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2055\,
            I => \N__2024\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2044\,
            I => \N__2015\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2033\,
            I => \N__2015\
        );

    \I__333\ : InMux
    port map (
            O => \N__2032\,
            I => \N__2010\
        );

    \I__332\ : InMux
    port map (
            O => \N__2031\,
            I => \N__2010\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__2024\,
            I => \N__2003\
        );

    \I__330\ : InMux
    port map (
            O => \N__2023\,
            I => \N__1994\
        );

    \I__329\ : InMux
    port map (
            O => \N__2022\,
            I => \N__1994\
        );

    \I__328\ : InMux
    port map (
            O => \N__2021\,
            I => \N__1994\
        );

    \I__327\ : InMux
    port map (
            O => \N__2020\,
            I => \N__1994\
        );

    \I__326\ : Span4Mux_v
    port map (
            O => \N__2015\,
            I => \N__1989\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2010\,
            I => \N__1989\
        );

    \I__324\ : InMux
    port map (
            O => \N__2009\,
            I => \N__1980\
        );

    \I__323\ : InMux
    port map (
            O => \N__2008\,
            I => \N__1980\
        );

    \I__322\ : InMux
    port map (
            O => \N__2007\,
            I => \N__1980\
        );

    \I__321\ : InMux
    port map (
            O => \N__2006\,
            I => \N__1980\
        );

    \I__320\ : Odrv4
    port map (
            O => \N__2003\,
            I => \S2_S3_c_1\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__1994\,
            I => \S2_S3_c_1\
        );

    \I__318\ : Odrv4
    port map (
            O => \N__1989\,
            I => \S2_S3_c_1\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1980\,
            I => \S2_S3_c_1\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__1971\,
            I => \SYNTHESIZED_WIRE_0_6_cascade_\
        );

    \I__315\ : InMux
    port map (
            O => \N__1968\,
            I => \N__1958\
        );

    \I__314\ : InMux
    port map (
            O => \N__1967\,
            I => \N__1955\
        );

    \I__313\ : InMux
    port map (
            O => \N__1966\,
            I => \N__1950\
        );

    \I__312\ : InMux
    port map (
            O => \N__1965\,
            I => \N__1950\
        );

    \I__311\ : InMux
    port map (
            O => \N__1964\,
            I => \N__1947\
        );

    \I__310\ : InMux
    port map (
            O => \N__1963\,
            I => \N__1942\
        );

    \I__309\ : InMux
    port map (
            O => \N__1962\,
            I => \N__1942\
        );

    \I__308\ : InMux
    port map (
            O => \N__1961\,
            I => \N__1939\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1958\,
            I => \N__1936\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1955\,
            I => \N__1929\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1950\,
            I => \N__1929\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1947\,
            I => \N__1929\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1942\,
            I => \N__1924\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1939\,
            I => \N__1924\
        );

    \I__301\ : Span4Mux_v
    port map (
            O => \N__1936\,
            I => \N__1919\
        );

    \I__300\ : Span4Mux_v
    port map (
            O => \N__1929\,
            I => \N__1919\
        );

    \I__299\ : Span4Mux_v
    port map (
            O => \N__1924\,
            I => \N__1916\
        );

    \I__298\ : Span4Mux_v
    port map (
            O => \N__1919\,
            I => \N__1913\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__1916\,
            I => \N__1910\
        );

    \I__296\ : Odrv4
    port map (
            O => \N__1913\,
            I => \S1_c\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__1910\,
            I => \S1_c\
        );

    \I__294\ : InMux
    port map (
            O => \N__1905\,
            I => \N__1902\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1902\,
            I => \b2v_inst4.result_reg2_bmZ0Z_6\
        );

    \I__292\ : InMux
    port map (
            O => \N__1899\,
            I => \N__1896\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1896\,
            I => \b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4\
        );

    \I__290\ : InMux
    port map (
            O => \N__1893\,
            I => \b2v_inst.un8_result_arith_cry_0\
        );

    \I__289\ : InMux
    port map (
            O => \N__1890\,
            I => \N__1887\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1887\,
            I => \b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4\
        );

    \I__287\ : InMux
    port map (
            O => \N__1884\,
            I => \b2v_inst.un8_result_arith_cry_1\
        );

    \I__286\ : InMux
    port map (
            O => \N__1881\,
            I => \N__1878\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1878\,
            I => \b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4\
        );

    \I__284\ : InMux
    port map (
            O => \N__1875\,
            I => \b2v_inst.un8_result_arith_cry_2\
        );

    \I__283\ : InMux
    port map (
            O => \N__1872\,
            I => \N__1869\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1869\,
            I => \un8_result_arith_cry_3_c_RNIO6R4\
        );

    \I__281\ : InMux
    port map (
            O => \N__1866\,
            I => \b2v_inst.un8_result_arith_cry_3\
        );

    \I__280\ : InMux
    port map (
            O => \N__1863\,
            I => \N__1860\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1860\,
            I => \b2v_inst3.result_reg1_amZ0Z_3\
        );

    \I__278\ : InMux
    port map (
            O => \N__1857\,
            I => \N__1854\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1854\,
            I => \b2v_inst.A_equal_B_NEZ0Z_1\
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__1851\,
            I => \b2v_inst3.result_reg1_bmZ0Z_2_cascade_\
        );

    \I__275\ : InMux
    port map (
            O => \N__1848\,
            I => \N__1845\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1845\,
            I => \b2v_inst3.result_reg1_amZ0Z_2\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__1842\,
            I => \SYNTHESIZED_WIRE_3_2_cascade_\
        );

    \I__272\ : IoInMux
    port map (
            O => \N__1839\,
            I => \N__1836\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1836\,
            I => \N__1833\
        );

    \I__270\ : Span4Mux_s0_h
    port map (
            O => \N__1833\,
            I => \N__1830\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__1830\,
            I => \N__1827\
        );

    \I__268\ : Odrv4
    port map (
            O => \N__1827\,
            I => \SYNTHESIZED_WIRE_4_2\
        );

    \I__267\ : InMux
    port map (
            O => \N__1824\,
            I => \N__1821\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1821\,
            I => \b2v_inst.A_equal_B_NEZ0Z_3\
        );

    \I__265\ : InMux
    port map (
            O => \N__1818\,
            I => \N__1815\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1815\,
            I => \b2v_inst.result_arith_1_2\
        );

    \I__263\ : InMux
    port map (
            O => \N__1812\,
            I => \N__1809\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1809\,
            I => \N_23\
        );

    \I__261\ : InMux
    port map (
            O => \N__1806\,
            I => \N__1794\
        );

    \I__260\ : InMux
    port map (
            O => \N__1805\,
            I => \N__1794\
        );

    \I__259\ : InMux
    port map (
            O => \N__1804\,
            I => \N__1789\
        );

    \I__258\ : InMux
    port map (
            O => \N__1803\,
            I => \N__1789\
        );

    \I__257\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1784\
        );

    \I__256\ : InMux
    port map (
            O => \N__1801\,
            I => \N__1784\
        );

    \I__255\ : InMux
    port map (
            O => \N__1800\,
            I => \N__1781\
        );

    \I__254\ : InMux
    port map (
            O => \N__1799\,
            I => \N__1778\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1794\,
            I => \N__1773\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__1789\,
            I => \N__1773\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1784\,
            I => \N__1770\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1781\,
            I => \N__1761\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1778\,
            I => \N__1761\
        );

    \I__248\ : Sp12to4
    port map (
            O => \N__1773\,
            I => \N__1761\
        );

    \I__247\ : Sp12to4
    port map (
            O => \N__1770\,
            I => \N__1761\
        );

    \I__246\ : Span12Mux_v
    port map (
            O => \N__1761\,
            I => \N__1758\
        );

    \I__245\ : Odrv12
    port map (
            O => \N__1758\,
            I => s2_c
        );

    \I__244\ : IoInMux
    port map (
            O => \N__1755\,
            I => \N__1752\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1752\,
            I => \N__1749\
        );

    \I__242\ : Odrv12
    port map (
            O => \N__1749\,
            I => \SYNTHESIZED_WIRE_4_6\
        );

    \I__241\ : InMux
    port map (
            O => \N__1746\,
            I => \N__1743\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1743\,
            I => \b2v_inst.A_c_i_6\
        );

    \I__239\ : InMux
    port map (
            O => \N__1740\,
            I => \N__1737\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1737\,
            I => \b2v_inst.A_c_i_7\
        );

    \I__237\ : InMux
    port map (
            O => \N__1734\,
            I => \bfn_1_14_0_\
        );

    \I__236\ : IoInMux
    port map (
            O => \N__1731\,
            I => \N__1727\
        );

    \I__235\ : CascadeMux
    port map (
            O => \N__1730\,
            I => \N__1724\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1727\,
            I => \N__1721\
        );

    \I__233\ : InMux
    port map (
            O => \N__1724\,
            I => \N__1718\
        );

    \I__232\ : Span4Mux_s2_v
    port map (
            O => \N__1721\,
            I => \N__1715\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1718\,
            I => \N__1712\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__1715\,
            I => \B_bigger_c_THRU_CO\
        );

    \I__229\ : Odrv4
    port map (
            O => \N__1712\,
            I => \B_bigger_c_THRU_CO\
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__1707\,
            I => \b2v_inst3.result_reg1_amZ0Z_1_cascade_\
        );

    \I__227\ : InMux
    port map (
            O => \N__1704\,
            I => \N__1701\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1701\,
            I => \b2v_inst3.result_reg1_bmZ0Z_1\
        );

    \I__225\ : InMux
    port map (
            O => \N__1698\,
            I => \N__1695\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1695\,
            I => \SYNTHESIZED_WIRE_3_1\
        );

    \I__223\ : CascadeMux
    port map (
            O => \N__1692\,
            I => \b2v_inst3.result_reg1_bmZ0Z_3_cascade_\
        );

    \I__222\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1686\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1686\,
            I => \SYNTHESIZED_WIRE_3_3\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__1683\,
            I => \N__1680\
        );

    \I__219\ : InMux
    port map (
            O => \N__1680\,
            I => \N__1677\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1677\,
            I => b2v_inst_result_arith_1_7
        );

    \I__217\ : InMux
    port map (
            O => \N__1674\,
            I => \b2v_inst.result_arith_1_cry_6\
        );

    \I__216\ : InMux
    port map (
            O => \N__1671\,
            I => \bfn_1_12_0_\
        );

    \I__215\ : IoInMux
    port map (
            O => \N__1668\,
            I => \N__1665\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1665\,
            I => \N__1662\
        );

    \I__213\ : IoSpan4Mux
    port map (
            O => \N__1662\,
            I => \N__1659\
        );

    \I__212\ : Sp12to4
    port map (
            O => \N__1659\,
            I => \N__1656\
        );

    \I__211\ : Span12Mux_s7_v
    port map (
            O => \N__1656\,
            I => \N__1653\
        );

    \I__210\ : Odrv12
    port map (
            O => \N__1653\,
            I => carry_out_c
        );

    \I__209\ : InMux
    port map (
            O => \N__1650\,
            I => \N__1647\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1647\,
            I => \b2v_inst.A_c_i_0\
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__1644\,
            I => \N__1641\
        );

    \I__206\ : InMux
    port map (
            O => \N__1641\,
            I => \N__1638\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1638\,
            I => \b2v_inst.A_c_i_1\
        );

    \I__204\ : CascadeMux
    port map (
            O => \N__1635\,
            I => \N__1632\
        );

    \I__203\ : InMux
    port map (
            O => \N__1632\,
            I => \N__1629\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1629\,
            I => \b2v_inst.A_c_i_2\
        );

    \I__201\ : InMux
    port map (
            O => \N__1626\,
            I => \N__1623\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1623\,
            I => \b2v_inst.A_c_i_3\
        );

    \I__199\ : InMux
    port map (
            O => \N__1620\,
            I => \N__1617\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1617\,
            I => \b2v_inst.A_c_i_4\
        );

    \I__197\ : InMux
    port map (
            O => \N__1614\,
            I => \N__1611\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1611\,
            I => \b2v_inst.A_c_i_5\
        );

    \I__195\ : CascadeMux
    port map (
            O => \N__1608\,
            I => \b2v_inst4.result_reg2_amZ0Z_7_cascade_\
        );

    \I__194\ : IoInMux
    port map (
            O => \N__1605\,
            I => \N__1602\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1602\,
            I => \SYNTHESIZED_WIRE_4_7\
        );

    \I__192\ : InMux
    port map (
            O => \N__1599\,
            I => \N__1596\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1596\,
            I => \b2v_inst.result_arith_1_1\
        );

    \I__190\ : InMux
    port map (
            O => \N__1593\,
            I => \b2v_inst.result_arith_1_cry_0\
        );

    \I__189\ : InMux
    port map (
            O => \N__1590\,
            I => \b2v_inst.result_arith_1_cry_1\
        );

    \I__188\ : InMux
    port map (
            O => \N__1587\,
            I => \N__1584\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1584\,
            I => \b2v_inst.result_arith_1_3\
        );

    \I__186\ : InMux
    port map (
            O => \N__1581\,
            I => \b2v_inst.result_arith_1_cry_2\
        );

    \I__185\ : CascadeMux
    port map (
            O => \N__1578\,
            I => \N__1575\
        );

    \I__184\ : InMux
    port map (
            O => \N__1575\,
            I => \N__1572\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1572\,
            I => b2v_inst_result_arith_1_4
        );

    \I__182\ : InMux
    port map (
            O => \N__1569\,
            I => \b2v_inst.result_arith_1_cry_3\
        );

    \I__181\ : CascadeMux
    port map (
            O => \N__1566\,
            I => \N__1563\
        );

    \I__180\ : InMux
    port map (
            O => \N__1563\,
            I => \N__1560\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1560\,
            I => b2v_inst_result_arith_1_5
        );

    \I__178\ : InMux
    port map (
            O => \N__1557\,
            I => \b2v_inst.result_arith_1_cry_4\
        );

    \I__177\ : InMux
    port map (
            O => \N__1554\,
            I => \b2v_inst.result_arith_1_cry_5\
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1551\,
            I => \b2v_inst4.result_reg2_bmZ0Z_4_cascade_\
        );

    \I__175\ : IoInMux
    port map (
            O => \N__1548\,
            I => \N__1545\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1545\,
            I => \N__1542\
        );

    \I__173\ : IoSpan4Mux
    port map (
            O => \N__1542\,
            I => \N__1539\
        );

    \I__172\ : Odrv4
    port map (
            O => \N__1539\,
            I => \SYNTHESIZED_WIRE_4_4\
        );

    \I__171\ : CascadeMux
    port map (
            O => \N__1536\,
            I => \SYNTHESIZED_WIRE_0_5_cascade_\
        );

    \I__170\ : CascadeMux
    port map (
            O => \N__1533\,
            I => \b2v_inst4.result_reg2_bmZ0Z_5_cascade_\
        );

    \I__169\ : IoInMux
    port map (
            O => \N__1530\,
            I => \N__1527\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1527\,
            I => \SYNTHESIZED_WIRE_4_5\
        );

    \I__167\ : CascadeMux
    port map (
            O => \N__1524\,
            I => \N__1521\
        );

    \I__166\ : InMux
    port map (
            O => \N__1521\,
            I => \N__1518\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1518\,
            I => \N__1515\
        );

    \I__164\ : Odrv12
    port map (
            O => \N__1515\,
            I => \N_22\
        );

    \I__163\ : CascadeMux
    port map (
            O => \N__1512\,
            I => \N_24_cascade_\
        );

    \I__162\ : IoInMux
    port map (
            O => \N__1509\,
            I => \N__1506\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1506\,
            I => \N__1503\
        );

    \I__160\ : Span4Mux_s0_h
    port map (
            O => \N__1503\,
            I => \N__1500\
        );

    \I__159\ : Span4Mux_v
    port map (
            O => \N__1500\,
            I => \N__1497\
        );

    \I__158\ : Odrv4
    port map (
            O => \N__1497\,
            I => \SYNTHESIZED_WIRE_4_3\
        );

    \I__157\ : InMux
    port map (
            O => \N__1494\,
            I => \N__1491\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1491\,
            I => \b2v_inst4.result_reg2_amZ0Z_4\
        );

    \I__155\ : InMux
    port map (
            O => \N__1488\,
            I => \N__1485\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1485\,
            I => \b2v_inst4.result_reg2_amZ0Z_5\
        );

    \I__153\ : IoInMux
    port map (
            O => \N__1482\,
            I => \N__1479\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1479\,
            I => \N__1476\
        );

    \I__151\ : Span4Mux_s0_h
    port map (
            O => \N__1476\,
            I => \N__1473\
        );

    \I__150\ : Odrv4
    port map (
            O => \N__1473\,
            I => \SYNTHESIZED_WIRE_4_1\
        );

    \I__149\ : InMux
    port map (
            O => \N__1470\,
            I => \N__1467\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1467\,
            I => \b2v_inst3.result_reg1_bmZ0Z_0\
        );

    \I__147\ : CascadeMux
    port map (
            O => \N__1464\,
            I => \b2v_inst3.result_reg1_amZ0Z_0_cascade_\
        );

    \I__146\ : CascadeMux
    port map (
            O => \N__1461\,
            I => \SYNTHESIZED_WIRE_3_0_cascade_\
        );

    \I__145\ : InMux
    port map (
            O => \N__1458\,
            I => \N__1455\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1455\,
            I => \N_21\
        );

    \I__143\ : IoInMux
    port map (
            O => \N__1452\,
            I => \N__1449\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1449\,
            I => \N__1446\
        );

    \I__141\ : IoSpan4Mux
    port map (
            O => \N__1446\,
            I => \N__1443\
        );

    \I__140\ : Odrv4
    port map (
            O => \N__1443\,
            I => \SYNTHESIZED_WIRE_4_0\
        );

    \I__139\ : CascadeMux
    port map (
            O => \N__1440\,
            I => \b2v_inst.A_equal_B_NEZ0Z_2_cascade_\
        );

    \I__138\ : InMux
    port map (
            O => \N__1437\,
            I => \N__1434\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1434\,
            I => \b2v_inst.A_equal_B_NEZ0Z_0\
        );

    \I__136\ : IoInMux
    port map (
            O => \N__1431\,
            I => \N__1428\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1428\,
            I => \N__1425\
        );

    \I__134\ : IoSpan4Mux
    port map (
            O => \N__1425\,
            I => \N__1422\
        );

    \I__133\ : IoSpan4Mux
    port map (
            O => \N__1422\,
            I => \N__1419\
        );

    \I__132\ : Odrv4
    port map (
            O => \N__1419\,
            I => \A_equal_B_c\
        );

    \I__131\ : CascadeMux
    port map (
            O => \N__1416\,
            I => \SYNTHESIZED_WIRE_0_4_cascade_\
        );

    \I__130\ : ClkMux
    port map (
            O => \N__1413\,
            I => \N__1398\
        );

    \I__129\ : ClkMux
    port map (
            O => \N__1412\,
            I => \N__1398\
        );

    \I__128\ : ClkMux
    port map (
            O => \N__1411\,
            I => \N__1398\
        );

    \I__127\ : ClkMux
    port map (
            O => \N__1410\,
            I => \N__1398\
        );

    \I__126\ : ClkMux
    port map (
            O => \N__1409\,
            I => \N__1398\
        );

    \I__125\ : GlobalMux
    port map (
            O => \N__1398\,
            I => \N__1395\
        );

    \I__124\ : gio2CtrlBuf
    port map (
            O => \N__1395\,
            I => \CLK_c_g\
        );

    \I__123\ : IoInMux
    port map (
            O => \N__1392\,
            I => \N__1389\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__1389\,
            I => \CONSTANT_ONE_NET\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.result_arith_1_8\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \B_bigger_c\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \A_bigger_c\,
            carryinitout => \bfn_2_13_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_bm_0_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__2322\,
            in1 => \N__2007\,
            in2 => \N__2146\,
            in3 => \N__2667\,
            lcout => \b2v_inst3.result_reg1_bmZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_0_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111010110100"
        )
    port map (
            in0 => \N__2120\,
            in1 => \N__2785\,
            in2 => \N__2844\,
            in3 => \N__2786\,
            lcout => \N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_equal_B_NE_0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__2577\,
            in1 => \N__2666\,
            in2 => \N__2843\,
            in3 => \N__2784\,
            lcout => \b2v_inst.A_equal_B_NEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_1_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__2009\,
            in1 => \N__1802\,
            in2 => \N__1524\,
            in3 => \N__1698\,
            lcout => \SYNTHESIZED_WIRE_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_am_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001100100"
        )
    port map (
            in0 => \N__2838\,
            in1 => \N__2006\,
            in2 => \N__2790\,
            in3 => \N__2121\,
            lcout => OPEN,
            ltout => \b2v_inst3.result_reg1_amZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_ns_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__1470\,
            in1 => \_gnd_net_\,
            in2 => \N__1464\,
            in3 => \N__1961\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__1801\,
            in1 => \N__2008\,
            in2 => \N__1461\,
            in3 => \N__1458\,
            lcout => \SYNTHESIZED_WIRE_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_equal_B_NE_2_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__3263\,
            in1 => \N__3217\,
            in2 => \N__3324\,
            in3 => \N__3379\,
            lcout => OPEN,
            ltout => \b2v_inst.A_equal_B_NEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_equal_B_NE_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1857\,
            in1 => \N__1824\,
            in2 => \N__1440\,
            in3 => \N__1437\,
            lcout => \A_equal_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.result_logic_4_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001100100"
        )
    port map (
            in0 => \N__3322\,
            in1 => \N__2020\,
            in2 => \N__2151\,
            in3 => \N__3380\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_bm_4_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__2022\,
            in1 => \N__1962\,
            in2 => \N__1416\,
            in3 => \N__2324\,
            lcout => OPEN,
            ltout => \b2v_inst4.result_reg2_bmZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_ns_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1803\,
            in2 => \N__1551\,
            in3 => \N__1494\,
            lcout => \SYNTHESIZED_WIRE_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.result_logic_5_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010011101010"
        )
    port map (
            in0 => \N__2021\,
            in1 => \N__2133\,
            in2 => \N__3225\,
            in3 => \N__3264\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_bm_5_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__1963\,
            in1 => \N__3381\,
            in2 => \N__1536\,
            in3 => \N__2023\,
            lcout => OPEN,
            ltout => \b2v_inst4.result_reg2_bmZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_ns_5_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__1804\,
            in1 => \_gnd_net_\,
            in2 => \N__1533\,
            in3 => \N__1488\,
            lcout => \SYNTHESIZED_WIRE_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_0_c_RNI1KOT_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__1599\,
            in1 => \N__1899\,
            in2 => \_gnd_net_\,
            in3 => \N__2186\,
            lcout => \N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_2_c_RNIB2TT_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2187\,
            in1 => \N__1881\,
            in2 => \_gnd_net_\,
            in3 => \N__1587\,
            lcout => OPEN,
            ltout => \N_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_3_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__1805\,
            in1 => \N__1689\,
            in2 => \N__1512\,
            in3 => \N__2080\,
            lcout => \SYNTHESIZED_WIRE_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_am_4_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__1872\,
            in1 => \N__2081\,
            in2 => \N__1578\,
            in3 => \N__2188\,
            lcout => \b2v_inst4.result_reg2_amZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_am_5_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__2189\,
            in1 => \N__2871\,
            in2 => \N__1566\,
            in3 => \N__2082\,
            lcout => \b2v_inst4.result_reg2_amZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_am_7_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__2083\,
            in1 => \N__2850\,
            in2 => \N__1683\,
            in3 => \N__2190\,
            lcout => OPEN,
            ltout => \b2v_inst4.result_reg2_amZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_ns_7_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__2220\,
            in1 => \_gnd_net_\,
            in2 => \N__1608\,
            in3 => \N__1806\,
            lcout => \SYNTHESIZED_WIRE_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_0_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2805\,
            in2 => \N__2782\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \b2v_inst.result_arith_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_0_c_RNIOBEO_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2549\,
            in2 => \N__2664\,
            in3 => \N__1593\,
            lcout => \b2v_inst.result_arith_1_1\,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_0\,
            carryout => \b2v_inst.result_arith_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_1_c_RNIRFFO_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2515\,
            in2 => \N__2436\,
            in3 => \N__1590\,
            lcout => \b2v_inst.result_arith_1_2\,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_1\,
            carryout => \b2v_inst.result_arith_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_2_c_RNIUJGO_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2379\,
            in2 => \N__2331\,
            in3 => \N__1581\,
            lcout => \b2v_inst.result_arith_1_3\,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_2\,
            carryout => \b2v_inst.result_arith_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_3_c_RNI1OHO_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3306\,
            in2 => \N__3378\,
            in3 => \N__1569\,
            lcout => b2v_inst_result_arith_1_4,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_3\,
            carryout => \b2v_inst.result_arith_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_4_c_RNI4SIO_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3252\,
            in2 => \N__3222\,
            in3 => \N__1557\,
            lcout => b2v_inst_result_arith_1_5,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_4\,
            carryout => \b2v_inst.result_arith_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_5_c_RNI70KO_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3124\,
            in2 => \N__3083\,
            in3 => \N__1554\,
            lcout => b2v_inst_result_arith_1_6,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_5\,
            carryout => \b2v_inst.result_arith_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_6_c_RNIA4LO_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2990\,
            in2 => \N__2947\,
            in3 => \N__1674\,
            lcout => b2v_inst_result_arith_1_7,
            ltout => OPEN,
            carryin => \b2v_inst.result_arith_1_cry_6\,
            carryout => \b2v_inst.result_arith_1_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.result_arith_1_cry_7_c_RNIQ27A_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__2191\,
            in1 => \N__2084\,
            in2 => \N__1730\,
            in3 => \N__1671\,
            lcout => carry_out_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_0_c_inv_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2751\,
            in1 => \N__1650\,
            in2 => \N__2842\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.A_c_i_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \b2v_inst.B_bigger_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_1_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2576\,
            in2 => \N__1644\,
            in3 => \N__2643\,
            lcout => \b2v_inst.A_c_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_0\,
            carryout => \b2v_inst.B_bigger_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_2_c_inv_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2501\,
            in1 => \N__2421\,
            in2 => \N__1635\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.A_c_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_1\,
            carryout => \b2v_inst.B_bigger_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_3_c_inv_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2287\,
            in1 => \N__1626\,
            in2 => \N__2378\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.A_c_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_2\,
            carryout => \b2v_inst.B_bigger_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_4_c_inv_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1620\,
            in2 => \N__3323\,
            in3 => \N__3340\,
            lcout => \b2v_inst.A_c_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_3\,
            carryout => \b2v_inst.B_bigger_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_5_c_inv_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3199\,
            in1 => \N__1614\,
            in2 => \N__3257\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.A_c_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_4\,
            carryout => \b2v_inst.B_bigger_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_6_c_inv_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3043\,
            in1 => \N__1746\,
            in2 => \N__3111\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.A_c_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_5\,
            carryout => \b2v_inst.B_bigger_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.B_bigger_cry_7_c_inv_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1740\,
            in2 => \N__3000\,
            in3 => \N__2910\,
            lcout => \b2v_inst.A_c_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.B_bigger_cry_6\,
            carryout => \B_bigger_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_bigger_c_THRU_LUT4_0_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1734\,
            lcout => \B_bigger_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_bm_1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__2771\,
            in1 => \N__2032\,
            in2 => \N__2516\,
            in3 => \N__2150\,
            lcout => \b2v_inst3.result_reg1_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_am_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010011101010"
        )
    port map (
            in0 => \N__2031\,
            in1 => \N__2657\,
            in2 => \N__2185\,
            in3 => \N__2575\,
            lcout => OPEN,
            ltout => \b2v_inst3.result_reg1_amZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_ns_1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__1964\,
            in1 => \_gnd_net_\,
            in2 => \N__1707\,
            in3 => \N__1704\,
            lcout => \SYNTHESIZED_WIRE_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_bm_3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__2195\,
            in1 => \N__2071\,
            in2 => \N__2783\,
            in3 => \N__2494\,
            lcout => OPEN,
            ltout => \b2v_inst3.result_reg1_bmZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_ns_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1863\,
            in2 => \N__1692\,
            in3 => \N__1966\,
            lcout => \SYNTHESIZED_WIRE_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_am_2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000101100"
        )
    port map (
            in0 => \N__2192\,
            in1 => \N__2068\,
            in2 => \N__2448\,
            in3 => \N__2493\,
            lcout => \b2v_inst3.result_reg1_amZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_am_3_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001001010"
        )
    port map (
            in0 => \N__2069\,
            in1 => \N__2193\,
            in2 => \N__2377\,
            in3 => \N__2329\,
            lcout => \b2v_inst3.result_reg1_amZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_equal_B_NE_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__2328\,
            in1 => \N__2367\,
            in2 => \N__2447\,
            in3 => \N__2492\,
            lcout => \b2v_inst.A_equal_B_NEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_bm_2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__2070\,
            in1 => \N__2330\,
            in2 => \N__2665\,
            in3 => \N__2194\,
            lcout => OPEN,
            ltout => \b2v_inst3.result_reg1_bmZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.result_reg1_ns_2_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__1965\,
            in1 => \_gnd_net_\,
            in2 => \N__1851\,
            in3 => \N__1848\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_2_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__2072\,
            in1 => \N__1812\,
            in2 => \N__1842\,
            in3 => \N__1799\,
            lcout => \SYNTHESIZED_WIRE_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_equal_B_NE_3_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3014\,
            in1 => \N__3125\,
            in2 => \N__3090\,
            in3 => \N__2948\,
            lcout => \b2v_inst.A_equal_B_NEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_1_c_RNI6RQT_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2196\,
            in1 => \N__1890\,
            in2 => \_gnd_net_\,
            in3 => \N__1818\,
            lcout => \N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_ns_6_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2208\,
            in1 => \N__1800\,
            in2 => \_gnd_net_\,
            in3 => \N__1905\,
            lcout => \SYNTHESIZED_WIRE_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.result_logic_7_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010011101010"
        )
    port map (
            in0 => \N__2074\,
            in1 => \N__2201\,
            in2 => \N__2952\,
            in3 => \N__3015\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_bm_7_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__3089\,
            in1 => \N__2079\,
            in2 => \N__2223\,
            in3 => \N__1968\,
            lcout => \b2v_inst4.result_reg2_bmZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_am_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__2197\,
            in1 => \N__2862\,
            in2 => \N__2085\,
            in3 => \N__2214\,
            lcout => \b2v_inst4.result_reg2_amZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.result_logic_6_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001011101100"
        )
    port map (
            in0 => \N__3088\,
            in1 => \N__2073\,
            in2 => \N__2202\,
            in3 => \N__3126\,
            lcout => OPEN,
            ltout => \SYNTHESIZED_WIRE_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.result_reg2_bm_6_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__2078\,
            in1 => \N__3223\,
            in2 => \N__1971\,
            in3 => \N__1967\,
            lcout => \b2v_inst4.result_reg2_bmZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_0_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2681\,
            in2 => \N__2770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \b2v_inst.un8_result_arith_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_0_c_RNIITN4_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2529\,
            in2 => \N__2663\,
            in3 => \N__1893\,
            lcout => \b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_0\,
            carryout => \b2v_inst.un8_result_arith_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_1_c_RNIK0P4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2391\,
            in2 => \N__2517\,
            in3 => \N__1884\,
            lcout => \b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_1\,
            carryout => \b2v_inst.un8_result_arith_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_2_c_RNIM3Q4_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2235\,
            in2 => \N__2323\,
            in3 => \N__1875\,
            lcout => \b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_2\,
            carryout => \b2v_inst.un8_result_arith_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_3_c_RNIO6R4_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3369\,
            in2 => \N__3279\,
            in3 => \N__1866\,
            lcout => \un8_result_arith_cry_3_c_RNIO6R4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_3\,
            carryout => \b2v_inst.un8_result_arith_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_4_c_RNIQ9S4_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3138\,
            in2 => \N__3221\,
            in3 => \N__2865\,
            lcout => \un8_result_arith_cry_4_c_RNIQ9S4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_4\,
            carryout => \b2v_inst.un8_result_arith_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_5_c_RNISCT4_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3027\,
            in2 => \N__3084\,
            in3 => \N__2856\,
            lcout => \un8_result_arith_cry_5_c_RNISCT4\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_result_arith_cry_5\,
            carryout => \b2v_inst.un8_result_arith_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_result_arith_cry_6_c_RNIK5GH_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__3012\,
            in1 => \N__2937\,
            in2 => \_gnd_net_\,
            in3 => \N__2853\,
            lcout => \un8_result_arith_cry_6_c_RNIK5GH\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_0_c_inv_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2831\,
            in1 => \N__2744\,
            in2 => \N__2682\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.B_c_i_0\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \b2v_inst.A_bigger_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_1_c_inv_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2528\,
            in2 => \N__2650\,
            in3 => \N__2574\,
            lcout => \b2v_inst.B_c_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_0\,
            carryout => \b2v_inst.A_bigger_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_2_c_inv_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2390\,
            in2 => \N__2511\,
            in3 => \N__2446\,
            lcout => \b2v_inst.B_c_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_1\,
            carryout => \b2v_inst.A_bigger_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_3_c_inv_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2360\,
            in1 => \N__2234\,
            in2 => \N__2311\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.B_c_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_2\,
            carryout => \b2v_inst.A_bigger_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_4_c_inv_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3275\,
            in2 => \N__3377\,
            in3 => \N__3307\,
            lcout => \b2v_inst.B_c_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_3\,
            carryout => \b2v_inst.A_bigger_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_5_c_inv_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3256\,
            in1 => \N__3137\,
            in2 => \N__3224\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.B_c_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_4\,
            carryout => \b2v_inst.A_bigger_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_6_c_inv_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3123\,
            in1 => \N__3026\,
            in2 => \N__3082\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.B_c_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_5\,
            carryout => \b2v_inst.A_bigger_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.A_bigger_cry_7_c_inv_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3013\,
            in1 => \N__2892\,
            in2 => \N__2946\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.B_c_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.A_bigger_cry_6\,
            carryout => \A_bigger_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \A_bigger_c_THRU_LUT4_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2886\,
            lcout => \A_bigger_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
