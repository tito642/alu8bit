-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 22 2023 21:20:02

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "alu_behavioral" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of alu_behavioral
entity alu_behavioral is
port (
    alu_out : out std_logic_vector(7 downto 0);
    s : in std_logic_vector(3 downto 0);
    A : in std_logic_vector(7 downto 0);
    B : in std_logic_vector(7 downto 0);
    clk : in std_logic);
end alu_behavioral;

-- Architecture of alu_behavioral
-- View name is \INTERFACE\
architecture \INTERFACE\ of alu_behavioral is

signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1837\ : std_logic;
signal \N__1834\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1755\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1621\ : std_logic;
signal \N__1618\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1581\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1539\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1468\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1450\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1417\ : std_logic;
signal \N__1414\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1405\ : std_logic;
signal \N__1404\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1392\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1384\ : std_logic;
signal \N__1381\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1375\ : std_logic;
signal \N__1372\ : std_logic;
signal \N__1369\ : std_logic;
signal \N__1366\ : std_logic;
signal \N__1363\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1354\ : std_logic;
signal \N__1351\ : std_logic;
signal \N__1348\ : std_logic;
signal \N__1345\ : std_logic;
signal \N__1342\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1336\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1330\ : std_logic;
signal \N__1327\ : std_logic;
signal \N__1324\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1309\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1303\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1297\ : std_logic;
signal \N__1296\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1285\ : std_logic;
signal \N__1282\ : std_logic;
signal \N__1279\ : std_logic;
signal \N__1276\ : std_logic;
signal \N__1271\ : std_logic;
signal \N__1268\ : std_logic;
signal \N__1267\ : std_logic;
signal \N__1264\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1258\ : std_logic;
signal \N__1255\ : std_logic;
signal \N__1246\ : std_logic;
signal \N__1243\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1237\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1231\ : std_logic;
signal \N__1228\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1224\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1222\ : std_logic;
signal \N__1221\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1204\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal clk_c_g : std_logic;
signal \alu_out_RNO_2Z0Z_1_cascade_\ : std_logic;
signal \N_143_cascade_\ : std_logic;
signal alu_out_13_1 : std_logic;
signal \alu_out38_cascade_\ : std_logic;
signal \un1_alu_out43_1_3_cascade_\ : std_logic;
signal un1_alu_out43_1_i : std_logic;
signal un1_alu_out43_1_2 : std_logic;
signal alu_out40_0 : std_logic;
signal \N_90_cascade_\ : std_logic;
signal \alu_out_RNO_3Z0Z_1\ : std_logic;
signal alu_out_13_5 : std_logic;
signal \N_87_cascade_\ : std_logic;
signal alu_out_13_4 : std_logic;
signal alu_out_13_0 : std_logic;
signal alu_out_13_6 : std_logic;
signal \s_c_i_1_cascade_\ : std_logic;
signal \N_88\ : std_logic;
signal \un1_A_1_cascade_\ : std_logic;
signal \B_c_0\ : std_logic;
signal \alu_out_RNO_2Z0Z_0_cascade_\ : std_logic;
signal \N_142\ : std_logic;
signal \alu_out_RNO_3Z0Z_0\ : std_logic;
signal \B_c_1\ : std_logic;
signal \N_85_cascade_\ : std_logic;
signal \B_c_4\ : std_logic;
signal \alu_out_RNO_3Z0Z_4\ : std_logic;
signal \alu_out_RNO_2Z0Z_4_cascade_\ : std_logic;
signal \N_146\ : std_logic;
signal \A_c_4\ : std_logic;
signal \alu_out_RNO_2Z0Z_5_cascade_\ : std_logic;
signal \alu_out_RNO_3Z0Z_5\ : std_logic;
signal \N_147\ : std_logic;
signal \alu_out_RNO_2Z0Z_3_cascade_\ : std_logic;
signal \alu_out_RNO_3Z0Z_3\ : std_logic;
signal \N_145_cascade_\ : std_logic;
signal alu_out_13_3 : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_1\ : std_logic;
signal \alu_out_RNO_3Z0Z_2_cascade_\ : std_logic;
signal \alu_out_RNO_2Z0Z_2\ : std_logic;
signal \N_144_cascade_\ : std_logic;
signal alu_out_13_2 : std_logic;
signal \s_ibuf_RNI1HJVZ0Z_0\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \un1_A_1\ : std_logic;
signal \B_ibuf_RNIE5VR2Z0Z_0\ : std_logic;
signal \alu_out_RNO_1Z0Z_0\ : std_logic;
signal \un1_A_1_cry_0_c_THRU_CO\ : std_logic;
signal \B_ibuf_RNIH05C1Z0Z_1\ : std_logic;
signal \B_ibuf_RNI08QF1Z0Z_1\ : std_logic;
signal \alu_out_RNO_1Z0Z_1\ : std_logic;
signal \un1_A_1_cry_0\ : std_logic;
signal \B_ibuf_RNI2AQF1Z0Z_2\ : std_logic;
signal \alu_out_RNO_1Z0Z_2\ : std_logic;
signal \un1_A_1_cry_1\ : std_logic;
signal \B_ibuf_RNIJ25C1Z0Z_3\ : std_logic;
signal \alu_out_RNO_1Z0Z_3\ : std_logic;
signal \un1_A_1_cry_2\ : std_logic;
signal \B_ibuf_RNIK35C1Z0Z_4\ : std_logic;
signal \B_ibuf_RNI6EQF1Z0Z_4\ : std_logic;
signal \alu_out_RNO_1Z0Z_4\ : std_logic;
signal \un1_A_1_cry_3\ : std_logic;
signal \B_ibuf_RNI8GQF1Z0Z_5\ : std_logic;
signal \alu_out_RNO_1Z0Z_5\ : std_logic;
signal \un1_A_1_cry_4\ : std_logic;
signal \B_ibuf_RNIM55C1Z0Z_6\ : std_logic;
signal \alu_out_RNO_1Z0Z_6\ : std_logic;
signal \un1_A_1_cry_5\ : std_logic;
signal \un1_A_1_cry_6\ : std_logic;
signal s_c_3 : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal alu_out_13_7 : std_logic;
signal \un1_A_1_axb_7\ : std_logic;
signal \alu_out_RNO_3Z0Z_7\ : std_logic;
signal \N_91\ : std_logic;
signal \B_ibuf_RNII15C1Z0Z_2\ : std_logic;
signal \B_c_2\ : std_logic;
signal \N_86\ : std_logic;
signal \B_c_5\ : std_logic;
signal \N_89_cascade_\ : std_logic;
signal \B_ibuf_RNIL45C1Z0Z_5\ : std_logic;
signal s_c_i_1 : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \alu_out_RNO_2Z0Z_6_cascade_\ : std_logic;
signal \alu_out_RNO_3Z0Z_6\ : std_logic;
signal \N_148\ : std_logic;
signal \B_c_3\ : std_logic;
signal \A_c_3\ : std_logic;
signal \B_ibuf_RNI4CQF1Z0Z_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \B_c_6\ : std_logic;
signal \B_ibuf_RNIAIQF1Z0Z_6\ : std_logic;
signal \A_c_7\ : std_logic;
signal s_c_1 : std_logic;
signal s_c_0 : std_logic;
signal \B_c_7\ : std_logic;
signal s_c_2 : std_logic;
signal \alu_out_RNO_5Z0Z_7\ : std_logic;
signal \alu_out_RNO_4Z0Z_7_cascade_\ : std_logic;
signal \N_149\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal \A_wire\ : std_logic_vector(7 downto 0);
signal \B_wire\ : std_logic_vector(7 downto 0);
signal alu_out_wire : std_logic_vector(7 downto 0);
signal s_wire : std_logic_vector(3 downto 0);

begin
    clk_wire <= clk;
    \A_wire\ <= A;
    \B_wire\ <= B;
    alu_out <= alu_out_wire;
    s_wire <= s;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2966\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2968\,
            DIN => \N__2967\,
            DOUT => \N__2966\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2968\,
            PADOUT => \N__2967\,
            PADIN => \N__2966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2957\,
            DIN => \N__2956\,
            DOUT => \N__2955\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2957\,
            PADOUT => \N__2956\,
            PADIN => \N__2955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2948\,
            DIN => \N__2947\,
            DOUT => \N__2946\,
            PACKAGEPIN => \B_wire\(7)
        );

    \B_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2948\,
            PADOUT => \N__2947\,
            PADIN => \N__2946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2939\,
            DIN => \N__2938\,
            DOUT => \N__2937\,
            PACKAGEPIN => alu_out_wire(6)
        );

    \alu_out_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2939\,
            PADOUT => \N__2938\,
            PADIN => \N__2937\,
            CLOCKENABLE => \N__1292\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1336\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1223\
        );

    \s_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2930\,
            DIN => \N__2929\,
            DOUT => \N__2928\,
            PACKAGEPIN => s_wire(0)
        );

    \s_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2930\,
            PADOUT => \N__2929\,
            PADIN => \N__2928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => s_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2921\,
            DIN => \N__2920\,
            DOUT => \N__2919\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2921\,
            PADOUT => \N__2920\,
            PADIN => \N__2919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2912\,
            DIN => \N__2911\,
            DOUT => \N__2910\,
            PACKAGEPIN => \B_wire\(3)
        );

    \B_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2912\,
            PADOUT => \N__2911\,
            PADIN => \N__2910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2903\,
            DIN => \N__2902\,
            DOUT => \N__2901\,
            PACKAGEPIN => alu_out_wire(3)
        );

    \alu_out_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2903\,
            PADOUT => \N__2902\,
            PADIN => \N__2901\,
            CLOCKENABLE => \N__1291\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1684\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1222\
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2894\,
            DIN => \N__2893\,
            DOUT => \N__2892\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2894\,
            PADOUT => \N__2893\,
            PADIN => \N__2892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2885\,
            DIN => \N__2884\,
            DOUT => \N__2883\,
            PACKAGEPIN => \B_wire\(6)
        );

    \B_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2885\,
            PADOUT => \N__2884\,
            PADIN => \N__2883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2876\,
            DIN => \N__2875\,
            DOUT => \N__2874\,
            PACKAGEPIN => alu_out_wire(7)
        );

    \alu_out_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2876\,
            PADOUT => \N__2875\,
            PADIN => \N__2874\,
            CLOCKENABLE => \N__1291\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1720\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1222\
        );

    \s_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2867\,
            DIN => \N__2866\,
            DOUT => \N__2865\,
            PACKAGEPIN => s_wire(1)
        );

    \s_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2867\,
            PADOUT => \N__2866\,
            PADIN => \N__2865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => s_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2858\,
            DIN => \N__2857\,
            DOUT => \N__2856\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2858\,
            PADOUT => \N__2857\,
            PADIN => \N__2856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2849\,
            DIN => \N__2848\,
            DOUT => \N__2847\,
            PACKAGEPIN => \B_wire\(2)
        );

    \B_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2849\,
            PADOUT => \N__2848\,
            PADIN => \N__2847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2840\,
            DIN => \N__2839\,
            DOUT => \N__2838\,
            PACKAGEPIN => alu_out_wire(0)
        );

    \alu_out_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2840\,
            PADOUT => \N__2839\,
            PADIN => \N__2838\,
            CLOCKENABLE => \N__1296\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1224\
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2831\,
            DIN => \N__2830\,
            DOUT => \N__2829\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2831\,
            PADOUT => \N__2830\,
            PADIN => \N__2829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2822\,
            DIN => \N__2821\,
            DOUT => \N__2820\,
            PACKAGEPIN => \B_wire\(0)
        );

    \B_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2822\,
            PADOUT => \N__2821\,
            PADIN => \N__2820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2813\,
            DIN => \N__2812\,
            DOUT => \N__2811\,
            PACKAGEPIN => alu_out_wire(2)
        );

    \alu_out_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2813\,
            PADOUT => \N__2812\,
            PADIN => \N__2811\,
            CLOCKENABLE => \N__1296\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1224\
        );

    \alu_out_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2804\,
            DIN => \N__2803\,
            DOUT => \N__2802\,
            PACKAGEPIN => alu_out_wire(4)
        );

    \alu_out_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2804\,
            PADOUT => \N__2803\,
            PADIN => \N__2802\,
            CLOCKENABLE => \N__1292\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1366\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1223\
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2795\,
            DIN => \N__2794\,
            DOUT => \N__2793\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2795\,
            PADOUT => \N__2794\,
            PADIN => \N__2793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2786\,
            DIN => \N__2785\,
            DOUT => \N__2784\,
            PACKAGEPIN => \B_wire\(5)
        );

    \B_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2786\,
            PADOUT => \N__2785\,
            PADIN => \N__2784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2777\,
            DIN => \N__2776\,
            DOUT => \N__2775\,
            PACKAGEPIN => alu_out_wire(1)
        );

    \alu_out_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2777\,
            PADOUT => \N__2776\,
            PADIN => \N__2775\,
            CLOCKENABLE => \N__1297\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1225\
        );

    \s_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2768\,
            DIN => \N__2767\,
            DOUT => \N__2766\,
            PACKAGEPIN => s_wire(2)
        );

    \s_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2768\,
            PADOUT => \N__2767\,
            PADIN => \N__2766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => s_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2759\,
            DIN => \N__2758\,
            DOUT => \N__2757\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2759\,
            PADOUT => \N__2758\,
            PADIN => \N__2757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2750\,
            DIN => \N__2749\,
            DOUT => \N__2748\,
            PACKAGEPIN => \B_wire\(1)
        );

    \B_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2750\,
            PADOUT => \N__2749\,
            PADIN => \N__2748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \alu_out_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2741\,
            DIN => \N__2740\,
            DOUT => \N__2739\,
            PACKAGEPIN => alu_out_wire(5)
        );

    \alu_out_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__2741\,
            PADOUT => \N__2740\,
            PADIN => \N__2739\,
            CLOCKENABLE => \N__1267\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1375\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1221\
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2732\,
            DIN => \N__2731\,
            DOUT => \N__2730\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2732\,
            PADOUT => \N__2731\,
            PADIN => \N__2730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2723\,
            DIN => \N__2722\,
            DOUT => \N__2721\,
            PACKAGEPIN => \B_wire\(4)
        );

    \B_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2723\,
            PADOUT => \N__2722\,
            PADIN => \N__2721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \B_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2714\,
            DIN => \N__2713\,
            DOUT => \N__2712\,
            PACKAGEPIN => s_wire(3)
        );

    \s_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2714\,
            PADOUT => \N__2713\,
            PADIN => \N__2712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => s_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__2695\,
            I => \alu_out_RNO_2Z0Z_6_cascade_\
        );

    \I__600\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__2689\,
            I => \alu_out_RNO_3Z0Z_6\
        );

    \I__598\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__2683\,
            I => \N__2680\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__2680\,
            I => \N_148\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__2677\,
            I => \N__2673\
        );

    \I__594\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2670\
        );

    \I__593\ : InMux
    port map (
            O => \N__2673\,
            I => \N__2666\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2670\,
            I => \N__2663\
        );

    \I__591\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2660\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__2666\,
            I => \N__2657\
        );

    \I__589\ : Span12Mux_s1_h
    port map (
            O => \N__2663\,
            I => \N__2652\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2660\,
            I => \N__2652\
        );

    \I__587\ : Odrv12
    port map (
            O => \N__2657\,
            I => \B_c_3\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__2652\,
            I => \B_c_3\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__2647\,
            I => \N__2644\
        );

    \I__584\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2637\
        );

    \I__583\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2637\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__2642\,
            I => \N__2634\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__2637\,
            I => \N__2630\
        );

    \I__580\ : InMux
    port map (
            O => \N__2634\,
            I => \N__2627\
        );

    \I__579\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2624\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__2630\,
            I => \N__2619\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2627\,
            I => \N__2619\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__2624\,
            I => \N__2616\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__2619\,
            I => \N__2613\
        );

    \I__574\ : Span4Mux_v
    port map (
            O => \N__2616\,
            I => \N__2610\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__2613\,
            I => \A_c_3\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__2610\,
            I => \A_c_3\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__570\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__2596\,
            I => \B_ibuf_RNI4CQF1Z0Z_3\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__2593\,
            I => \N__2588\
        );

    \I__566\ : InMux
    port map (
            O => \N__2592\,
            I => \N__2581\
        );

    \I__565\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2581\
        );

    \I__564\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2581\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__2581\,
            I => \N__2577\
        );

    \I__562\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2574\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__2577\,
            I => \A_c_6\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2574\,
            I => \A_c_6\
        );

    \I__559\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2564\
        );

    \I__558\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2559\
        );

    \I__557\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2559\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__2564\,
            I => \N__2556\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2559\,
            I => \N__2553\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__2556\,
            I => \N__2550\
        );

    \I__553\ : Span12Mux_s5_v
    port map (
            O => \N__2553\,
            I => \N__2547\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__2550\,
            I => \B_c_6\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__2547\,
            I => \B_c_6\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__2542\,
            I => \N__2539\
        );

    \I__549\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2536\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2536\,
            I => \N__2533\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__2533\,
            I => \B_ibuf_RNIAIQF1Z0Z_6\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__2530\,
            I => \N__2525\
        );

    \I__545\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2520\
        );

    \I__544\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2520\
        );

    \I__543\ : InMux
    port map (
            O => \N__2525\,
            I => \N__2517\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__2520\,
            I => \N__2514\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2517\,
            I => \N__2510\
        );

    \I__540\ : Span4Mux_h
    port map (
            O => \N__2514\,
            I => \N__2507\
        );

    \I__539\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2504\
        );

    \I__538\ : Span12Mux_s11_h
    port map (
            O => \N__2510\,
            I => \N__2501\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__2507\,
            I => \N__2498\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2504\,
            I => \N__2495\
        );

    \I__535\ : Odrv12
    port map (
            O => \N__2501\,
            I => \A_c_7\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__2498\,
            I => \A_c_7\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__2495\,
            I => \A_c_7\
        );

    \I__532\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2469\
        );

    \I__531\ : InMux
    port map (
            O => \N__2487\,
            I => \N__2469\
        );

    \I__530\ : InMux
    port map (
            O => \N__2486\,
            I => \N__2469\
        );

    \I__529\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2469\
        );

    \I__528\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2466\
        );

    \I__527\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2459\
        );

    \I__526\ : InMux
    port map (
            O => \N__2482\,
            I => \N__2459\
        );

    \I__525\ : InMux
    port map (
            O => \N__2481\,
            I => \N__2459\
        );

    \I__524\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2452\
        );

    \I__523\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2452\
        );

    \I__522\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2452\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2469\,
            I => \N__2446\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__2466\,
            I => \N__2446\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2459\,
            I => \N__2441\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__2452\,
            I => \N__2441\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__2451\,
            I => \N__2434\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__2446\,
            I => \N__2428\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__2441\,
            I => \N__2425\
        );

    \I__514\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2418\
        );

    \I__513\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2418\
        );

    \I__512\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2418\
        );

    \I__511\ : InMux
    port map (
            O => \N__2437\,
            I => \N__2411\
        );

    \I__510\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2411\
        );

    \I__509\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2411\
        );

    \I__508\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2406\
        );

    \I__507\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2406\
        );

    \I__506\ : Sp12to4
    port map (
            O => \N__2428\,
            I => \N__2399\
        );

    \I__505\ : Sp12to4
    port map (
            O => \N__2425\,
            I => \N__2399\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2418\,
            I => \N__2399\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2411\,
            I => s_c_1
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2406\,
            I => s_c_1
        );

    \I__501\ : Odrv12
    port map (
            O => \N__2399\,
            I => s_c_1
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__2392\,
            I => \N__2386\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__2391\,
            I => \N__2383\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__2390\,
            I => \N__2368\
        );

    \I__497\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2352\
        );

    \I__496\ : InMux
    port map (
            O => \N__2386\,
            I => \N__2352\
        );

    \I__495\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2352\
        );

    \I__494\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2352\
        );

    \I__493\ : InMux
    port map (
            O => \N__2381\,
            I => \N__2347\
        );

    \I__492\ : InMux
    port map (
            O => \N__2380\,
            I => \N__2347\
        );

    \I__491\ : InMux
    port map (
            O => \N__2379\,
            I => \N__2338\
        );

    \I__490\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2338\
        );

    \I__489\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2338\
        );

    \I__488\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2338\
        );

    \I__487\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2327\
        );

    \I__486\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2327\
        );

    \I__485\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2327\
        );

    \I__484\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2327\
        );

    \I__483\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2327\
        );

    \I__482\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2318\
        );

    \I__481\ : InMux
    port map (
            O => \N__2367\,
            I => \N__2318\
        );

    \I__480\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2318\
        );

    \I__479\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2318\
        );

    \I__478\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2309\
        );

    \I__477\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2309\
        );

    \I__476\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2309\
        );

    \I__475\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2309\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2352\,
            I => \N__2304\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2347\,
            I => \N__2297\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2338\,
            I => \N__2297\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2297\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2318\,
            I => \N__2292\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2309\,
            I => \N__2292\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2308\,
            I => \N__2280\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__2307\,
            I => \N__2275\
        );

    \I__466\ : Span4Mux_v
    port map (
            O => \N__2304\,
            I => \N__2268\
        );

    \I__465\ : Span4Mux_v
    port map (
            O => \N__2297\,
            I => \N__2268\
        );

    \I__464\ : Span4Mux_v
    port map (
            O => \N__2292\,
            I => \N__2268\
        );

    \I__463\ : InMux
    port map (
            O => \N__2291\,
            I => \N__2259\
        );

    \I__462\ : InMux
    port map (
            O => \N__2290\,
            I => \N__2259\
        );

    \I__461\ : InMux
    port map (
            O => \N__2289\,
            I => \N__2259\
        );

    \I__460\ : InMux
    port map (
            O => \N__2288\,
            I => \N__2259\
        );

    \I__459\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2246\
        );

    \I__458\ : InMux
    port map (
            O => \N__2286\,
            I => \N__2246\
        );

    \I__457\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2246\
        );

    \I__456\ : InMux
    port map (
            O => \N__2284\,
            I => \N__2246\
        );

    \I__455\ : InMux
    port map (
            O => \N__2283\,
            I => \N__2246\
        );

    \I__454\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2246\
        );

    \I__453\ : InMux
    port map (
            O => \N__2279\,
            I => \N__2239\
        );

    \I__452\ : InMux
    port map (
            O => \N__2278\,
            I => \N__2239\
        );

    \I__451\ : InMux
    port map (
            O => \N__2275\,
            I => \N__2239\
        );

    \I__450\ : Odrv4
    port map (
            O => \N__2268\,
            I => s_c_0
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2259\,
            I => s_c_0
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2246\,
            I => s_c_0
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2239\,
            I => s_c_0
        );

    \I__446\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2225\
        );

    \I__445\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2222\
        );

    \I__444\ : InMux
    port map (
            O => \N__2228\,
            I => \N__2219\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2225\,
            I => \N__2216\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2222\,
            I => \N__2211\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2219\,
            I => \N__2211\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__2216\,
            I => \N__2208\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__2211\,
            I => \B_c_7\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__2208\,
            I => \B_c_7\
        );

    \I__437\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2192\
        );

    \I__436\ : InMux
    port map (
            O => \N__2202\,
            I => \N__2192\
        );

    \I__435\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2189\
        );

    \I__434\ : InMux
    port map (
            O => \N__2200\,
            I => \N__2184\
        );

    \I__433\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2184\
        );

    \I__432\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2179\
        );

    \I__431\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2179\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2192\,
            I => \N__2174\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2189\,
            I => \N__2174\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2184\,
            I => \N__2169\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2179\,
            I => \N__2169\
        );

    \I__426\ : Span4Mux_v
    port map (
            O => \N__2174\,
            I => \N__2162\
        );

    \I__425\ : Span4Mux_v
    port map (
            O => \N__2169\,
            I => \N__2159\
        );

    \I__424\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2150\
        );

    \I__423\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2150\
        );

    \I__422\ : InMux
    port map (
            O => \N__2166\,
            I => \N__2150\
        );

    \I__421\ : InMux
    port map (
            O => \N__2165\,
            I => \N__2150\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2162\,
            I => s_c_2
        );

    \I__419\ : Odrv4
    port map (
            O => \N__2159\,
            I => s_c_2
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2150\,
            I => s_c_2
        );

    \I__417\ : InMux
    port map (
            O => \N__2143\,
            I => \N__2140\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2140\,
            I => \alu_out_RNO_5Z0Z_7\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__2137\,
            I => \alu_out_RNO_4Z0Z_7_cascade_\
        );

    \I__414\ : InMux
    port map (
            O => \N__2134\,
            I => \N__2131\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2131\,
            I => \N_149\
        );

    \I__412\ : InMux
    port map (
            O => \N__2128\,
            I => \N__2125\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2125\,
            I => \alu_out_RNO_3Z0Z_7\
        );

    \I__410\ : InMux
    port map (
            O => \N__2122\,
            I => \N__2119\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2119\,
            I => \N_91\
        );

    \I__408\ : InMux
    port map (
            O => \N__2116\,
            I => \N__2113\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__2110\,
            I => \B_ibuf_RNII15C1Z0Z_2\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__2107\,
            I => \N__2103\
        );

    \I__404\ : InMux
    port map (
            O => \N__2106\,
            I => \N__2098\
        );

    \I__403\ : InMux
    port map (
            O => \N__2103\,
            I => \N__2098\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2098\,
            I => \N__2094\
        );

    \I__401\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2091\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__2094\,
            I => \N__2086\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2091\,
            I => \N__2086\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__2086\,
            I => \N__2083\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__2083\,
            I => \B_c_2\
        );

    \I__396\ : InMux
    port map (
            O => \N__2080\,
            I => \N__2077\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2077\,
            I => \N_86\
        );

    \I__394\ : InMux
    port map (
            O => \N__2074\,
            I => \N__2071\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2071\,
            I => \N__2067\
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__2070\,
            I => \N__2064\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__2067\,
            I => \N__2060\
        );

    \I__390\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2055\
        );

    \I__389\ : InMux
    port map (
            O => \N__2063\,
            I => \N__2055\
        );

    \I__388\ : Odrv4
    port map (
            O => \N__2060\,
            I => \B_c_5\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2055\,
            I => \B_c_5\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__2050\,
            I => \N_89_cascade_\
        );

    \I__385\ : InMux
    port map (
            O => \N__2047\,
            I => \N__2044\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2044\,
            I => \B_ibuf_RNIL45C1Z0Z_5\
        );

    \I__383\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2035\
        );

    \I__382\ : InMux
    port map (
            O => \N__2040\,
            I => \N__2027\
        );

    \I__381\ : InMux
    port map (
            O => \N__2039\,
            I => \N__2027\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__2038\,
            I => \N__2022\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2035\,
            I => \N__2016\
        );

    \I__378\ : InMux
    port map (
            O => \N__2034\,
            I => \N__2009\
        );

    \I__377\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2009\
        );

    \I__376\ : InMux
    port map (
            O => \N__2032\,
            I => \N__2009\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2027\,
            I => \N__2006\
        );

    \I__374\ : InMux
    port map (
            O => \N__2026\,
            I => \N__2001\
        );

    \I__373\ : InMux
    port map (
            O => \N__2025\,
            I => \N__2001\
        );

    \I__372\ : InMux
    port map (
            O => \N__2022\,
            I => \N__1994\
        );

    \I__371\ : InMux
    port map (
            O => \N__2021\,
            I => \N__1994\
        );

    \I__370\ : InMux
    port map (
            O => \N__2020\,
            I => \N__1994\
        );

    \I__369\ : InMux
    port map (
            O => \N__2019\,
            I => \N__1991\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__2016\,
            I => s_c_i_1
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2009\,
            I => s_c_i_1
        );

    \I__366\ : Odrv4
    port map (
            O => \N__2006\,
            I => s_c_i_1
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2001\,
            I => s_c_i_1
        );

    \I__364\ : LocalMux
    port map (
            O => \N__1994\,
            I => s_c_i_1
        );

    \I__363\ : LocalMux
    port map (
            O => \N__1991\,
            I => s_c_i_1
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__1978\,
            I => \N__1975\
        );

    \I__361\ : InMux
    port map (
            O => \N__1975\,
            I => \N__1971\
        );

    \I__360\ : InMux
    port map (
            O => \N__1974\,
            I => \N__1968\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__1971\,
            I => \N__1965\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__1968\,
            I => \N__1962\
        );

    \I__357\ : Span4Mux_v
    port map (
            O => \N__1965\,
            I => \N__1957\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__1962\,
            I => \N__1954\
        );

    \I__355\ : InMux
    port map (
            O => \N__1961\,
            I => \N__1949\
        );

    \I__354\ : InMux
    port map (
            O => \N__1960\,
            I => \N__1949\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__1957\,
            I => \A_c_0\
        );

    \I__352\ : Odrv4
    port map (
            O => \N__1954\,
            I => \A_c_0\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__1949\,
            I => \A_c_0\
        );

    \I__350\ : InMux
    port map (
            O => \N__1942\,
            I => \N__1939\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1939\,
            I => \N__1935\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__1938\,
            I => \N__1930\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__1935\,
            I => \N__1927\
        );

    \I__346\ : InMux
    port map (
            O => \N__1934\,
            I => \N__1924\
        );

    \I__345\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1919\
        );

    \I__344\ : InMux
    port map (
            O => \N__1930\,
            I => \N__1919\
        );

    \I__343\ : Odrv4
    port map (
            O => \N__1927\,
            I => \A_c_5\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1924\,
            I => \A_c_5\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__1919\,
            I => \A_c_5\
        );

    \I__340\ : InMux
    port map (
            O => \N__1912\,
            I => \N__1909\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__1909\,
            I => \B_ibuf_RNIH05C1Z0Z_1\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__1906\,
            I => \N__1903\
        );

    \I__337\ : InMux
    port map (
            O => \N__1903\,
            I => \N__1900\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1900\,
            I => \B_ibuf_RNI08QF1Z0Z_1\
        );

    \I__335\ : InMux
    port map (
            O => \N__1897\,
            I => \N__1894\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__1894\,
            I => \N__1891\
        );

    \I__333\ : Odrv4
    port map (
            O => \N__1891\,
            I => \alu_out_RNO_1Z0Z_1\
        );

    \I__332\ : InMux
    port map (
            O => \N__1888\,
            I => \un1_A_1_cry_0\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__1885\,
            I => \N__1882\
        );

    \I__330\ : InMux
    port map (
            O => \N__1882\,
            I => \N__1879\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__1879\,
            I => \B_ibuf_RNI2AQF1Z0Z_2\
        );

    \I__328\ : InMux
    port map (
            O => \N__1876\,
            I => \N__1873\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__1873\,
            I => \alu_out_RNO_1Z0Z_2\
        );

    \I__326\ : InMux
    port map (
            O => \N__1870\,
            I => \un1_A_1_cry_1\
        );

    \I__325\ : InMux
    port map (
            O => \N__1867\,
            I => \N__1864\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1864\,
            I => \B_ibuf_RNIJ25C1Z0Z_3\
        );

    \I__323\ : InMux
    port map (
            O => \N__1861\,
            I => \N__1858\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__1858\,
            I => \alu_out_RNO_1Z0Z_3\
        );

    \I__321\ : InMux
    port map (
            O => \N__1855\,
            I => \un1_A_1_cry_2\
        );

    \I__320\ : InMux
    port map (
            O => \N__1852\,
            I => \N__1849\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__1849\,
            I => \B_ibuf_RNIK35C1Z0Z_4\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__1846\,
            I => \N__1843\
        );

    \I__317\ : InMux
    port map (
            O => \N__1843\,
            I => \N__1840\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1840\,
            I => \B_ibuf_RNI6EQF1Z0Z_4\
        );

    \I__315\ : InMux
    port map (
            O => \N__1837\,
            I => \N__1834\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__1834\,
            I => \alu_out_RNO_1Z0Z_4\
        );

    \I__313\ : InMux
    port map (
            O => \N__1831\,
            I => \un1_A_1_cry_3\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__1828\,
            I => \N__1825\
        );

    \I__311\ : InMux
    port map (
            O => \N__1825\,
            I => \N__1822\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1822\,
            I => \N__1819\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__1819\,
            I => \B_ibuf_RNI8GQF1Z0Z_5\
        );

    \I__308\ : InMux
    port map (
            O => \N__1816\,
            I => \N__1813\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1813\,
            I => \alu_out_RNO_1Z0Z_5\
        );

    \I__306\ : InMux
    port map (
            O => \N__1810\,
            I => \un1_A_1_cry_4\
        );

    \I__305\ : InMux
    port map (
            O => \N__1807\,
            I => \N__1804\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1804\,
            I => \N__1801\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__1801\,
            I => \B_ibuf_RNIM55C1Z0Z_6\
        );

    \I__302\ : InMux
    port map (
            O => \N__1798\,
            I => \N__1795\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1795\,
            I => \alu_out_RNO_1Z0Z_6\
        );

    \I__300\ : InMux
    port map (
            O => \N__1792\,
            I => \un1_A_1_cry_5\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__1789\,
            I => \N__1786\
        );

    \I__298\ : InMux
    port map (
            O => \N__1786\,
            I => \N__1783\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1783\,
            I => \N__1774\
        );

    \I__296\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1769\
        );

    \I__295\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1769\
        );

    \I__294\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1760\
        );

    \I__293\ : InMux
    port map (
            O => \N__1779\,
            I => \N__1760\
        );

    \I__292\ : InMux
    port map (
            O => \N__1778\,
            I => \N__1760\
        );

    \I__291\ : InMux
    port map (
            O => \N__1777\,
            I => \N__1760\
        );

    \I__290\ : Span4Mux_v
    port map (
            O => \N__1774\,
            I => \N__1755\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__1769\,
            I => \N__1755\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1760\,
            I => \N__1752\
        );

    \I__287\ : Span4Mux_v
    port map (
            O => \N__1755\,
            I => \N__1745\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__1752\,
            I => \N__1742\
        );

    \I__285\ : InMux
    port map (
            O => \N__1751\,
            I => \N__1739\
        );

    \I__284\ : InMux
    port map (
            O => \N__1750\,
            I => \N__1732\
        );

    \I__283\ : InMux
    port map (
            O => \N__1749\,
            I => \N__1732\
        );

    \I__282\ : InMux
    port map (
            O => \N__1748\,
            I => \N__1732\
        );

    \I__281\ : Odrv4
    port map (
            O => \N__1745\,
            I => s_c_3
        );

    \I__280\ : Odrv4
    port map (
            O => \N__1742\,
            I => s_c_3
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1739\,
            I => s_c_3
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1732\,
            I => s_c_3
        );

    \I__277\ : InMux
    port map (
            O => \N__1723\,
            I => \bfn_2_11_0_\
        );

    \I__276\ : IoInMux
    port map (
            O => \N__1720\,
            I => \N__1717\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1717\,
            I => \N__1714\
        );

    \I__274\ : IoSpan4Mux
    port map (
            O => \N__1714\,
            I => \N__1711\
        );

    \I__273\ : Span4Mux_s1_h
    port map (
            O => \N__1711\,
            I => \N__1708\
        );

    \I__272\ : Span4Mux_h
    port map (
            O => \N__1708\,
            I => \N__1705\
        );

    \I__271\ : Odrv4
    port map (
            O => \N__1705\,
            I => alu_out_13_7
        );

    \I__270\ : InMux
    port map (
            O => \N__1702\,
            I => \N__1699\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1699\,
            I => \un1_A_1_axb_7\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__1696\,
            I => \alu_out_RNO_2Z0Z_3_cascade_\
        );

    \I__267\ : InMux
    port map (
            O => \N__1693\,
            I => \N__1690\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1690\,
            I => \alu_out_RNO_3Z0Z_3\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__1687\,
            I => \N_145_cascade_\
        );

    \I__264\ : IoInMux
    port map (
            O => \N__1684\,
            I => \N__1681\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1681\,
            I => \N__1678\
        );

    \I__262\ : Span4Mux_s2_h
    port map (
            O => \N__1678\,
            I => \N__1675\
        );

    \I__261\ : Odrv4
    port map (
            O => \N__1675\,
            I => alu_out_13_3
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1672\,
            I => \N__1669\
        );

    \I__259\ : InMux
    port map (
            O => \N__1669\,
            I => \N__1661\
        );

    \I__258\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1661\
        );

    \I__257\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1656\
        );

    \I__256\ : InMux
    port map (
            O => \N__1666\,
            I => \N__1656\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1661\,
            I => \N__1651\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1656\,
            I => \N__1651\
        );

    \I__253\ : Span4Mux_v
    port map (
            O => \N__1651\,
            I => \N__1648\
        );

    \I__252\ : Span4Mux_v
    port map (
            O => \N__1648\,
            I => \N__1645\
        );

    \I__251\ : Odrv4
    port map (
            O => \N__1645\,
            I => \A_c_2\
        );

    \I__250\ : InMux
    port map (
            O => \N__1642\,
            I => \N__1634\
        );

    \I__249\ : InMux
    port map (
            O => \N__1641\,
            I => \N__1634\
        );

    \I__248\ : InMux
    port map (
            O => \N__1640\,
            I => \N__1631\
        );

    \I__247\ : InMux
    port map (
            O => \N__1639\,
            I => \N__1628\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1634\,
            I => \N__1621\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1631\,
            I => \N__1621\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1628\,
            I => \N__1621\
        );

    \I__243\ : Span4Mux_v
    port map (
            O => \N__1621\,
            I => \N__1618\
        );

    \I__242\ : Span4Mux_v
    port map (
            O => \N__1618\,
            I => \N__1615\
        );

    \I__241\ : Odrv4
    port map (
            O => \N__1615\,
            I => \A_c_1\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__1612\,
            I => \alu_out_RNO_3Z0Z_2_cascade_\
        );

    \I__239\ : InMux
    port map (
            O => \N__1609\,
            I => \N__1606\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1606\,
            I => \alu_out_RNO_2Z0Z_2\
        );

    \I__237\ : CascadeMux
    port map (
            O => \N__1603\,
            I => \N_144_cascade_\
        );

    \I__236\ : IoInMux
    port map (
            O => \N__1600\,
            I => \N__1597\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1597\,
            I => \N__1594\
        );

    \I__234\ : Span12Mux_s1_h
    port map (
            O => \N__1594\,
            I => \N__1591\
        );

    \I__233\ : Odrv12
    port map (
            O => \N__1591\,
            I => alu_out_13_2
        );

    \I__232\ : CascadeMux
    port map (
            O => \N__1588\,
            I => \N__1585\
        );

    \I__231\ : InMux
    port map (
            O => \N__1585\,
            I => \N__1581\
        );

    \I__230\ : InMux
    port map (
            O => \N__1584\,
            I => \N__1578\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__1581\,
            I => \s_ibuf_RNI1HJVZ0Z_0\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1578\,
            I => \s_ibuf_RNI1HJVZ0Z_0\
        );

    \I__227\ : InMux
    port map (
            O => \N__1573\,
            I => \N__1570\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1570\,
            I => \un1_A_1\
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__1567\,
            I => \N__1564\
        );

    \I__224\ : InMux
    port map (
            O => \N__1564\,
            I => \N__1561\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1561\,
            I => \B_ibuf_RNIE5VR2Z0Z_0\
        );

    \I__222\ : InMux
    port map (
            O => \N__1558\,
            I => \N__1555\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1555\,
            I => \alu_out_RNO_1Z0Z_0\
        );

    \I__220\ : InMux
    port map (
            O => \N__1552\,
            I => \un1_A_1_cry_0_c_THRU_CO\
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__1549\,
            I => \N_85_cascade_\
        );

    \I__218\ : InMux
    port map (
            O => \N__1546\,
            I => \N__1540\
        );

    \I__217\ : InMux
    port map (
            O => \N__1545\,
            I => \N__1540\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1540\,
            I => \N__1536\
        );

    \I__215\ : CascadeMux
    port map (
            O => \N__1539\,
            I => \N__1533\
        );

    \I__214\ : Span4Mux_v
    port map (
            O => \N__1536\,
            I => \N__1530\
        );

    \I__213\ : InMux
    port map (
            O => \N__1533\,
            I => \N__1527\
        );

    \I__212\ : Odrv4
    port map (
            O => \N__1530\,
            I => \B_c_4\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1527\,
            I => \B_c_4\
        );

    \I__210\ : InMux
    port map (
            O => \N__1522\,
            I => \N__1519\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1519\,
            I => \alu_out_RNO_3Z0Z_4\
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__1516\,
            I => \alu_out_RNO_2Z0Z_4_cascade_\
        );

    \I__207\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1510\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1510\,
            I => \N__1507\
        );

    \I__205\ : Odrv4
    port map (
            O => \N__1507\,
            I => \N_146\
        );

    \I__204\ : InMux
    port map (
            O => \N__1504\,
            I => \N__1500\
        );

    \I__203\ : InMux
    port map (
            O => \N__1503\,
            I => \N__1497\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1500\,
            I => \N__1492\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1497\,
            I => \N__1489\
        );

    \I__200\ : InMux
    port map (
            O => \N__1496\,
            I => \N__1484\
        );

    \I__199\ : InMux
    port map (
            O => \N__1495\,
            I => \N__1484\
        );

    \I__198\ : Span4Mux_v
    port map (
            O => \N__1492\,
            I => \N__1477\
        );

    \I__197\ : Span4Mux_h
    port map (
            O => \N__1489\,
            I => \N__1477\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1484\,
            I => \N__1477\
        );

    \I__195\ : Span4Mux_v
    port map (
            O => \N__1477\,
            I => \N__1474\
        );

    \I__194\ : Odrv4
    port map (
            O => \N__1474\,
            I => \A_c_4\
        );

    \I__193\ : CascadeMux
    port map (
            O => \N__1471\,
            I => \alu_out_RNO_2Z0Z_5_cascade_\
        );

    \I__192\ : InMux
    port map (
            O => \N__1468\,
            I => \N__1465\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1465\,
            I => \alu_out_RNO_3Z0Z_5\
        );

    \I__190\ : InMux
    port map (
            O => \N__1462\,
            I => \N__1459\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1459\,
            I => \N__1456\
        );

    \I__188\ : Odrv12
    port map (
            O => \N__1456\,
            I => \N_147\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__1453\,
            I => \s_c_i_1_cascade_\
        );

    \I__186\ : InMux
    port map (
            O => \N__1450\,
            I => \N__1447\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1447\,
            I => \N_88\
        );

    \I__184\ : CascadeMux
    port map (
            O => \N__1444\,
            I => \un1_A_1_cascade_\
        );

    \I__183\ : CascadeMux
    port map (
            O => \N__1441\,
            I => \N__1437\
        );

    \I__182\ : CascadeMux
    port map (
            O => \N__1440\,
            I => \N__1434\
        );

    \I__181\ : InMux
    port map (
            O => \N__1437\,
            I => \N__1426\
        );

    \I__180\ : InMux
    port map (
            O => \N__1434\,
            I => \N__1426\
        );

    \I__179\ : InMux
    port map (
            O => \N__1433\,
            I => \N__1426\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1426\,
            I => \N__1423\
        );

    \I__177\ : Odrv12
    port map (
            O => \N__1423\,
            I => \B_c_0\
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1420\,
            I => \alu_out_RNO_2Z0Z_0_cascade_\
        );

    \I__175\ : InMux
    port map (
            O => \N__1417\,
            I => \N__1414\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1414\,
            I => \N_142\
        );

    \I__173\ : InMux
    port map (
            O => \N__1411\,
            I => \N__1408\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1408\,
            I => \alu_out_RNO_3Z0Z_0\
        );

    \I__171\ : InMux
    port map (
            O => \N__1405\,
            I => \N__1398\
        );

    \I__170\ : InMux
    port map (
            O => \N__1404\,
            I => \N__1398\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__1403\,
            I => \N__1395\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1398\,
            I => \N__1392\
        );

    \I__167\ : InMux
    port map (
            O => \N__1395\,
            I => \N__1389\
        );

    \I__166\ : Span4Mux_v
    port map (
            O => \N__1392\,
            I => \N__1384\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1389\,
            I => \N__1384\
        );

    \I__164\ : Span4Mux_v
    port map (
            O => \N__1384\,
            I => \N__1381\
        );

    \I__163\ : Span4Mux_v
    port map (
            O => \N__1381\,
            I => \N__1378\
        );

    \I__162\ : Odrv4
    port map (
            O => \N__1378\,
            I => \B_c_1\
        );

    \I__161\ : IoInMux
    port map (
            O => \N__1375\,
            I => \N__1372\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1372\,
            I => alu_out_13_5
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__1369\,
            I => \N_87_cascade_\
        );

    \I__158\ : IoInMux
    port map (
            O => \N__1366\,
            I => \N__1363\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1363\,
            I => \N__1360\
        );

    \I__156\ : IoSpan4Mux
    port map (
            O => \N__1360\,
            I => \N__1357\
        );

    \I__155\ : Span4Mux_s0_h
    port map (
            O => \N__1357\,
            I => \N__1354\
        );

    \I__154\ : Odrv4
    port map (
            O => \N__1354\,
            I => alu_out_13_4
        );

    \I__153\ : IoInMux
    port map (
            O => \N__1351\,
            I => \N__1348\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1348\,
            I => \N__1345\
        );

    \I__151\ : IoSpan4Mux
    port map (
            O => \N__1345\,
            I => \N__1342\
        );

    \I__150\ : Span4Mux_s0_h
    port map (
            O => \N__1342\,
            I => \N__1339\
        );

    \I__149\ : Odrv4
    port map (
            O => \N__1339\,
            I => alu_out_13_0
        );

    \I__148\ : IoInMux
    port map (
            O => \N__1336\,
            I => \N__1333\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1333\,
            I => \N__1330\
        );

    \I__146\ : Span4Mux_s0_h
    port map (
            O => \N__1330\,
            I => \N__1327\
        );

    \I__145\ : Span4Mux_v
    port map (
            O => \N__1327\,
            I => \N__1324\
        );

    \I__144\ : Odrv4
    port map (
            O => \N__1324\,
            I => alu_out_13_6
        );

    \I__143\ : CascadeMux
    port map (
            O => \N__1321\,
            I => \N_143_cascade_\
        );

    \I__142\ : IoInMux
    port map (
            O => \N__1318\,
            I => \N__1315\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1315\,
            I => \N__1312\
        );

    \I__140\ : Span4Mux_s0_h
    port map (
            O => \N__1312\,
            I => \N__1309\
        );

    \I__139\ : Span4Mux_v
    port map (
            O => \N__1309\,
            I => \N__1306\
        );

    \I__138\ : Odrv4
    port map (
            O => \N__1306\,
            I => alu_out_13_1
        );

    \I__137\ : CascadeMux
    port map (
            O => \N__1303\,
            I => \alu_out38_cascade_\
        );

    \I__136\ : CascadeMux
    port map (
            O => \N__1300\,
            I => \un1_alu_out43_1_3_cascade_\
        );

    \I__135\ : CEMux
    port map (
            O => \N__1297\,
            I => \N__1293\
        );

    \I__134\ : CEMux
    port map (
            O => \N__1296\,
            I => \N__1288\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1293\,
            I => \N__1285\
        );

    \I__132\ : CEMux
    port map (
            O => \N__1292\,
            I => \N__1282\
        );

    \I__131\ : CEMux
    port map (
            O => \N__1291\,
            I => \N__1279\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1288\,
            I => \N__1276\
        );

    \I__129\ : IoSpan4Mux
    port map (
            O => \N__1285\,
            I => \N__1271\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__1282\,
            I => \N__1271\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1279\,
            I => \N__1268\
        );

    \I__126\ : Span4Mux_s1_h
    port map (
            O => \N__1276\,
            I => \N__1264\
        );

    \I__125\ : IoSpan4Mux
    port map (
            O => \N__1271\,
            I => \N__1261\
        );

    \I__124\ : Span4Mux_s0_h
    port map (
            O => \N__1268\,
            I => \N__1258\
        );

    \I__123\ : CEMux
    port map (
            O => \N__1267\,
            I => \N__1255\
        );

    \I__122\ : Odrv4
    port map (
            O => \N__1264\,
            I => un1_alu_out43_1_i
        );

    \I__121\ : Odrv4
    port map (
            O => \N__1261\,
            I => un1_alu_out43_1_i
        );

    \I__120\ : Odrv4
    port map (
            O => \N__1258\,
            I => un1_alu_out43_1_i
        );

    \I__119\ : LocalMux
    port map (
            O => \N__1255\,
            I => un1_alu_out43_1_i
        );

    \I__118\ : InMux
    port map (
            O => \N__1246\,
            I => \N__1243\
        );

    \I__117\ : LocalMux
    port map (
            O => \N__1243\,
            I => un1_alu_out43_1_2
        );

    \I__116\ : InMux
    port map (
            O => \N__1240\,
            I => \N__1237\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__1237\,
            I => alu_out40_0
        );

    \I__114\ : CascadeMux
    port map (
            O => \N__1234\,
            I => \N_90_cascade_\
        );

    \I__113\ : InMux
    port map (
            O => \N__1231\,
            I => \N__1228\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1228\,
            I => \alu_out_RNO_3Z0Z_1\
        );

    \I__111\ : ClkMux
    port map (
            O => \N__1225\,
            I => \N__1210\
        );

    \I__110\ : ClkMux
    port map (
            O => \N__1224\,
            I => \N__1210\
        );

    \I__109\ : ClkMux
    port map (
            O => \N__1223\,
            I => \N__1210\
        );

    \I__108\ : ClkMux
    port map (
            O => \N__1222\,
            I => \N__1210\
        );

    \I__107\ : ClkMux
    port map (
            O => \N__1221\,
            I => \N__1210\
        );

    \I__106\ : GlobalMux
    port map (
            O => \N__1210\,
            I => \N__1207\
        );

    \I__105\ : gio2CtrlBuf
    port map (
            O => \N__1207\,
            I => clk_c_g
        );

    \I__104\ : CascadeMux
    port map (
            O => \N__1204\,
            I => \alu_out_RNO_2Z0Z_1_cascade_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_A_1_cry_6\,
            carryinitout => \bfn_2_11_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \alu_out_RNO_2_1_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001101000"
        )
    port map (
            in0 => \N__2365\,
            in1 => \N__2433\,
            in2 => \N__1403\,
            in3 => \N__1639\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_1_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2165\,
            in1 => \_gnd_net_\,
            in2 => \N__1204\,
            in3 => \N__1231\,
            lcout => OPEN,
            ltout => \N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__1777\,
            in1 => \_gnd_net_\,
            in2 => \N__1321\,
            in3 => \N__1897\,
            lcout => alu_out_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNI667V1_0_2_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2166\,
            in1 => \N__1779\,
            in2 => \N__2451\,
            in3 => \N__2367\,
            lcout => OPEN,
            ltout => \alu_out38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNID58E4_2_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__1240\,
            in1 => \N__2040\,
            in2 => \N__1303\,
            in3 => \N__2168\,
            lcout => OPEN,
            ltout => \un1_alu_out43_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNIJBFD6_2_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1300\,
            in3 => \N__1246\,
            lcout => un1_alu_out43_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNI667V1_2_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101110111"
        )
    port map (
            in0 => \N__1780\,
            in1 => \N__2167\,
            in2 => \N__2390\,
            in3 => \N__2437\,
            lcout => un1_alu_out43_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNI4CDF1_3_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__2039\,
            in1 => \N__1778\,
            in2 => \_gnd_net_\,
            in3 => \N__2366\,
            lcout => alu_out40_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNILCBS_6_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2289\,
            in2 => \_gnd_net_\,
            in3 => \N__2569\,
            lcout => OPEN,
            ltout => \N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIM55C1_6_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1234\,
            in3 => \N__2026\,
            lcout => \B_ibuf_RNIM55C1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_1_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__1974\,
            in1 => \N__1666\,
            in2 => \_gnd_net_\,
            in3 => \N__2290\,
            lcout => \alu_out_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_5_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__1751\,
            in1 => \N__1816\,
            in2 => \_gnd_net_\,
            in3 => \N__1462\,
            lcout => alu_out_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNII9BS_3_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2676\,
            in2 => \_gnd_net_\,
            in3 => \N__2288\,
            lcout => OPEN,
            ltout => \N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIJ25C1_3_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1369\,
            in3 => \N__2025\,
            lcout => \B_ibuf_RNIJ25C1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_3_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__1504\,
            in1 => \N__2291\,
            in2 => \_gnd_net_\,
            in3 => \N__1667\,
            lcout => \alu_out_RNO_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_4_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__1749\,
            in1 => \N__1837\,
            in2 => \_gnd_net_\,
            in3 => \N__1513\,
            lcout => alu_out_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNI6EQF1_4_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__2431\,
            in1 => \N__1545\,
            in2 => \N__2307\,
            in3 => \N__1503\,
            lcout => \B_ibuf_RNI6EQF1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIJABS_4_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__1546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2278\,
            lcout => \N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__1558\,
            in1 => \N__1748\,
            in2 => \_gnd_net_\,
            in3 => \N__1417\,
            lcout => alu_out_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNI1HJV_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2279\,
            lcout => \s_ibuf_RNI1HJVZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_6_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__1798\,
            in1 => \N__1750\,
            in2 => \_gnd_net_\,
            in3 => \N__2686\,
            lcout => alu_out_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \s_ibuf_RNI1PPF_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2432\,
            lcout => s_c_i_1,
            ltout => \s_c_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIK35C1_4_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1453\,
            in3 => \N__1450\,
            lcout => \B_ibuf_RNIK35C1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNI08QF1_1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__1641\,
            in1 => \N__2478\,
            in2 => \N__2308\,
            in3 => \N__1404\,
            lcout => \B_ibuf_RNI08QF1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIU5QF1_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__2479\,
            in1 => \N__2285\,
            in2 => \N__1440\,
            in3 => \N__1960\,
            lcout => \un1_A_1\,
            ltout => \un1_A_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIE5VR2_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__2283\,
            in1 => \N__2020\,
            in2 => \N__1444\,
            in3 => \N__1433\,
            lcout => \B_ibuf_RNIE5VR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111001101000"
        )
    port map (
            in0 => \N__2480\,
            in1 => \N__2286\,
            in2 => \N__1441\,
            in3 => \N__1961\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2201\,
            in2 => \N__1420\,
            in3 => \N__1411\,
            lcout => \N_142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_0_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__2513\,
            in1 => \N__1642\,
            in2 => \N__2038\,
            in3 => \N__2287\,
            lcout => \alu_out_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIG7BS_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1405\,
            lcout => OPEN,
            ltout => \N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIH05C1_1_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__2021\,
            in1 => \_gnd_net_\,
            in2 => \N__1549\,
            in3 => \_gnd_net_\,
            lcout => \B_ibuf_RNIH05C1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_4_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2633\,
            in1 => \N__2374\,
            in2 => \_gnd_net_\,
            in3 => \N__1934\,
            lcout => \alu_out_RNO_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_4_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001101000"
        )
    port map (
            in0 => \N__2372\,
            in1 => \N__2482\,
            in2 => \N__1539\,
            in3 => \N__1495\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_4_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__1522\,
            in1 => \_gnd_net_\,
            in2 => \N__1516\,
            in3 => \N__2202\,
            lcout => \N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_5_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2375\,
            in1 => \N__2580\,
            in2 => \_gnd_net_\,
            in3 => \N__1496\,
            lcout => \alu_out_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNI8GQF1_5_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__2481\,
            in1 => \N__2063\,
            in2 => \N__1938\,
            in3 => \N__2371\,
            lcout => \B_ibuf_RNI8GQF1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_5_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001101000"
        )
    port map (
            in0 => \N__2373\,
            in1 => \N__2483\,
            in2 => \N__2070\,
            in3 => \N__1933\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_5_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2203\,
            in2 => \N__1471\,
            in3 => \N__1468\,
            lcout => \N_147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111001101000"
        )
    port map (
            in0 => \N__2440\,
            in1 => \N__2363\,
            in2 => \N__2677\,
            in3 => \N__2643\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2198\,
            in1 => \_gnd_net_\,
            in2 => \N__1696\,
            in3 => \N__1693\,
            lcout => OPEN,
            ltout => \N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__1861\,
            in1 => \_gnd_net_\,
            in2 => \N__1687\,
            in3 => \N__1782\,
            lcout => alu_out_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNI2AQF1_2_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__2361\,
            in1 => \N__2438\,
            in2 => \N__2107\,
            in3 => \N__1668\,
            lcout => \B_ibuf_RNI2AQF1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_2_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011101000"
        )
    port map (
            in0 => \N__2439\,
            in1 => \N__2362\,
            in2 => \N__1672\,
            in3 => \N__2106\,
            lcout => \alu_out_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2364\,
            in1 => \_gnd_net_\,
            in2 => \N__2647\,
            in3 => \N__1640\,
            lcout => OPEN,
            ltout => \alu_out_RNO_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_2_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2197\,
            in2 => \N__1612\,
            in3 => \N__1609\,
            lcout => OPEN,
            ltout => \N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__1781\,
            in1 => \_gnd_net_\,
            in2 => \N__1603\,
            in3 => \N__1876\,
            lcout => alu_out_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_A_1_cry_0_c_THRU_CRY_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1584\,
            in2 => \N__1588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \un1_A_1_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1573\,
            in2 => \N__1567\,
            in3 => \N__1552\,
            lcout => \alu_out_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_0_c_THRU_CO\,
            carryout => \un1_A_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1912\,
            in2 => \N__1906\,
            in3 => \N__1888\,
            lcout => \alu_out_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_0\,
            carryout => \un1_A_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2116\,
            in2 => \N__1885\,
            in3 => \N__1870\,
            lcout => \alu_out_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_1\,
            carryout => \un1_A_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_3_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1867\,
            in2 => \N__2605\,
            in3 => \N__1855\,
            lcout => \alu_out_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_2\,
            carryout => \un1_A_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_4_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1852\,
            in2 => \N__1846\,
            in3 => \N__1831\,
            lcout => \alu_out_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_3\,
            carryout => \un1_A_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_5_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2047\,
            in2 => \N__1828\,
            in3 => \N__1810\,
            lcout => \alu_out_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_4\,
            carryout => \un1_A_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_6_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1807\,
            in2 => \N__2542\,
            in3 => \N__1792\,
            lcout => \alu_out_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \un1_A_1_cry_5\,
            carryout => \un1_A_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_7_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__2134\,
            in1 => \N__1702\,
            in2 => \N__1789\,
            in3 => \N__1723\,
            lcout => alu_out_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_7_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__2122\,
            in1 => \N__2034\,
            in2 => \_gnd_net_\,
            in3 => \N__2128\,
            lcout => \un1_A_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_7_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__2484\,
            in1 => \N__2379\,
            in2 => \N__2530\,
            in3 => \N__2229\,
            lcout => \alu_out_RNO_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_7_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2228\,
            lcout => \N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNII15C1_2_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2080\,
            lcout => \B_ibuf_RNII15C1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIH8BS_2_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2097\,
            lcout => \N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIKBBS_5_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2377\,
            lcout => OPEN,
            ltout => \N_89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIL45C1_5_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2050\,
            in3 => \N__2033\,
            lcout => \B_ibuf_RNIL45C1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_5_7_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__2389\,
            in1 => \N__2041\,
            in2 => \N__1978\,
            in3 => \N__2592\,
            lcout => \alu_out_RNO_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_3_6_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2381\,
            in1 => \N__2528\,
            in2 => \_gnd_net_\,
            in3 => \N__1942\,
            lcout => \alu_out_RNO_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_2_6_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001101000"
        )
    port map (
            in0 => \N__2568\,
            in1 => \N__2487\,
            in2 => \N__2391\,
            in3 => \N__2591\,
            lcout => OPEN,
            ltout => \alu_out_RNO_2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_0_6_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2199\,
            in1 => \_gnd_net_\,
            in2 => \N__2695\,
            in3 => \N__2692\,
            lcout => \N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNI4CQF1_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__2669\,
            in1 => \N__2485\,
            in2 => \N__2642\,
            in3 => \N__2380\,
            lcout => \B_ibuf_RNI4CQF1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \B_ibuf_RNIAIQF1_6_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__2486\,
            in1 => \N__2382\,
            in2 => \N__2593\,
            in3 => \N__2567\,
            lcout => \B_ibuf_RNIAIQF1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_4_7_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__2529\,
            in1 => \N__2488\,
            in2 => \N__2392\,
            in3 => \N__2230\,
            lcout => OPEN,
            ltout => \alu_out_RNO_4Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alu_out_RNO_1_7_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__2200\,
            in1 => \N__2143\,
            in2 => \N__2137\,
            in3 => \_gnd_net_\,
            lcout => \N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
