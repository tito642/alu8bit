// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 20 2023 04:45:29

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "ALU_STURCTURE" view "INTERFACE"

module ALU_STURCTURE (
    S2_S3,
    A,
    F,
    B,
    flag_zero,
    A_equal_B,
    B_bigger,
    s2,
    over_flow,
    carry_out,
    S1,
    A_bigger,
    CLK);

    input [1:0] S2_S3;
    input [7:0] A;
    output [7:0] F;
    input [7:0] B;
    output flag_zero;
    output A_equal_B;
    output B_bigger;
    input s2;
    output over_flow;
    output carry_out;
    input S1;
    output A_bigger;
    input CLK;

    wire N__3708;
    wire N__3707;
    wire N__3706;
    wire N__3697;
    wire N__3696;
    wire N__3695;
    wire N__3688;
    wire N__3687;
    wire N__3686;
    wire N__3679;
    wire N__3678;
    wire N__3677;
    wire N__3670;
    wire N__3669;
    wire N__3668;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3652;
    wire N__3651;
    wire N__3650;
    wire N__3643;
    wire N__3642;
    wire N__3641;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3625;
    wire N__3624;
    wire N__3623;
    wire N__3616;
    wire N__3615;
    wire N__3614;
    wire N__3607;
    wire N__3606;
    wire N__3605;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3589;
    wire N__3588;
    wire N__3587;
    wire N__3580;
    wire N__3579;
    wire N__3578;
    wire N__3571;
    wire N__3570;
    wire N__3569;
    wire N__3562;
    wire N__3561;
    wire N__3560;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3544;
    wire N__3543;
    wire N__3542;
    wire N__3535;
    wire N__3534;
    wire N__3533;
    wire N__3526;
    wire N__3525;
    wire N__3524;
    wire N__3517;
    wire N__3516;
    wire N__3515;
    wire N__3508;
    wire N__3507;
    wire N__3506;
    wire N__3499;
    wire N__3498;
    wire N__3497;
    wire N__3490;
    wire N__3489;
    wire N__3488;
    wire N__3481;
    wire N__3480;
    wire N__3479;
    wire N__3472;
    wire N__3471;
    wire N__3470;
    wire N__3463;
    wire N__3462;
    wire N__3461;
    wire N__3454;
    wire N__3453;
    wire N__3452;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3436;
    wire N__3435;
    wire N__3434;
    wire N__3427;
    wire N__3426;
    wire N__3425;
    wire N__3418;
    wire N__3417;
    wire N__3416;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3400;
    wire N__3399;
    wire N__3398;
    wire N__3381;
    wire N__3380;
    wire N__3379;
    wire N__3378;
    wire N__3377;
    wire N__3370;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3344;
    wire N__3341;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3324;
    wire N__3323;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3311;
    wire N__3308;
    wire N__3307;
    wire N__3306;
    wire N__3303;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3289;
    wire N__3286;
    wire N__3279;
    wire N__3276;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3264;
    wire N__3263;
    wire N__3258;
    wire N__3257;
    wire N__3256;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3225;
    wire N__3224;
    wire N__3223;
    wire N__3222;
    wire N__3221;
    wire N__3218;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3200;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3150;
    wire N__3147;
    wire N__3138;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3126;
    wire N__3125;
    wire N__3124;
    wire N__3123;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3111;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3090;
    wire N__3089;
    wire N__3088;
    wire N__3085;
    wire N__3084;
    wire N__3083;
    wire N__3082;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3047;
    wire N__3044;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3027;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3015;
    wire N__3014;
    wire N__3013;
    wire N__3012;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2959;
    wire N__2952;
    wire N__2949;
    wire N__2948;
    wire N__2947;
    wire N__2946;
    wire N__2941;
    wire N__2938;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2910;
    wire N__2907;
    wire N__2902;
    wire N__2899;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2843;
    wire N__2842;
    wire N__2839;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2831;
    wire N__2828;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2806;
    wire N__2805;
    wire N__2798;
    wire N__2795;
    wire N__2790;
    wire N__2787;
    wire N__2786;
    wire N__2785;
    wire N__2784;
    wire N__2783;
    wire N__2782;
    wire N__2775;
    wire N__2772;
    wire N__2771;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2715;
    wire N__2710;
    wire N__2707;
    wire N__2700;
    wire N__2697;
    wire N__2692;
    wire N__2689;
    wire N__2682;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2667;
    wire N__2666;
    wire N__2665;
    wire N__2664;
    wire N__2663;
    wire N__2658;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2595;
    wire N__2592;
    wire N__2587;
    wire N__2584;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2565;
    wire N__2562;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2549;
    wire N__2544;
    wire N__2539;
    wire N__2536;
    wire N__2529;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2517;
    wire N__2516;
    wire N__2515;
    wire N__2512;
    wire N__2511;
    wire N__2508;
    wire N__2505;
    wire N__2502;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2494;
    wire N__2493;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2470;
    wire N__2461;
    wire N__2456;
    wire N__2453;
    wire N__2448;
    wire N__2447;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2436;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2422;
    wire N__2421;
    wire N__2418;
    wire N__2415;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2398;
    wire N__2391;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2374;
    wire N__2371;
    wire N__2368;
    wire N__2367;
    wire N__2364;
    wire N__2361;
    wire N__2360;
    wire N__2355;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2331;
    wire N__2330;
    wire N__2329;
    wire N__2328;
    wire N__2325;
    wire N__2324;
    wire N__2323;
    wire N__2322;
    wire N__2315;
    wire N__2312;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2262;
    wire N__2259;
    wire N__2256;
    wire N__2251;
    wire N__2248;
    wire N__2245;
    wire N__2242;
    wire N__2235;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2211;
    wire N__2208;
    wire N__2205;
    wire N__2202;
    wire N__2201;
    wire N__2198;
    wire N__2197;
    wire N__2196;
    wire N__2195;
    wire N__2194;
    wire N__2193;
    wire N__2192;
    wire N__2191;
    wire N__2190;
    wire N__2189;
    wire N__2188;
    wire N__2187;
    wire N__2186;
    wire N__2185;
    wire N__2180;
    wire N__2175;
    wire N__2166;
    wire N__2163;
    wire N__2152;
    wire N__2151;
    wire N__2150;
    wire N__2147;
    wire N__2146;
    wire N__2139;
    wire N__2134;
    wire N__2133;
    wire N__2130;
    wire N__2125;
    wire N__2122;
    wire N__2121;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2109;
    wire N__2106;
    wire N__2103;
    wire N__2098;
    wire N__2085;
    wire N__2084;
    wire N__2083;
    wire N__2082;
    wire N__2081;
    wire N__2080;
    wire N__2079;
    wire N__2078;
    wire N__2075;
    wire N__2074;
    wire N__2073;
    wire N__2072;
    wire N__2071;
    wire N__2070;
    wire N__2069;
    wire N__2068;
    wire N__2065;
    wire N__2060;
    wire N__2055;
    wire N__2044;
    wire N__2033;
    wire N__2032;
    wire N__2031;
    wire N__2024;
    wire N__2023;
    wire N__2022;
    wire N__2021;
    wire N__2020;
    wire N__2015;
    wire N__2010;
    wire N__2009;
    wire N__2008;
    wire N__2007;
    wire N__2006;
    wire N__2003;
    wire N__1994;
    wire N__1989;
    wire N__1980;
    wire N__1971;
    wire N__1968;
    wire N__1967;
    wire N__1966;
    wire N__1965;
    wire N__1964;
    wire N__1963;
    wire N__1962;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1950;
    wire N__1947;
    wire N__1942;
    wire N__1939;
    wire N__1936;
    wire N__1929;
    wire N__1924;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1905;
    wire N__1902;
    wire N__1899;
    wire N__1896;
    wire N__1893;
    wire N__1890;
    wire N__1887;
    wire N__1884;
    wire N__1881;
    wire N__1878;
    wire N__1875;
    wire N__1872;
    wire N__1869;
    wire N__1866;
    wire N__1863;
    wire N__1860;
    wire N__1857;
    wire N__1854;
    wire N__1851;
    wire N__1848;
    wire N__1845;
    wire N__1842;
    wire N__1839;
    wire N__1836;
    wire N__1833;
    wire N__1830;
    wire N__1827;
    wire N__1824;
    wire N__1821;
    wire N__1818;
    wire N__1815;
    wire N__1812;
    wire N__1809;
    wire N__1806;
    wire N__1805;
    wire N__1804;
    wire N__1803;
    wire N__1802;
    wire N__1801;
    wire N__1800;
    wire N__1799;
    wire N__1794;
    wire N__1789;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1773;
    wire N__1770;
    wire N__1761;
    wire N__1758;
    wire N__1755;
    wire N__1752;
    wire N__1749;
    wire N__1746;
    wire N__1743;
    wire N__1740;
    wire N__1737;
    wire N__1734;
    wire N__1731;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1707;
    wire N__1704;
    wire N__1701;
    wire N__1698;
    wire N__1695;
    wire N__1692;
    wire N__1689;
    wire N__1686;
    wire N__1683;
    wire N__1680;
    wire N__1677;
    wire N__1674;
    wire N__1671;
    wire N__1668;
    wire N__1665;
    wire N__1662;
    wire N__1659;
    wire N__1656;
    wire N__1653;
    wire N__1650;
    wire N__1647;
    wire N__1644;
    wire N__1641;
    wire N__1638;
    wire N__1635;
    wire N__1632;
    wire N__1629;
    wire N__1626;
    wire N__1623;
    wire N__1620;
    wire N__1617;
    wire N__1614;
    wire N__1611;
    wire N__1608;
    wire N__1605;
    wire N__1602;
    wire N__1599;
    wire N__1596;
    wire N__1593;
    wire N__1590;
    wire N__1587;
    wire N__1584;
    wire N__1581;
    wire N__1578;
    wire N__1575;
    wire N__1572;
    wire N__1569;
    wire N__1566;
    wire N__1563;
    wire N__1560;
    wire N__1557;
    wire N__1554;
    wire N__1551;
    wire N__1548;
    wire N__1545;
    wire N__1542;
    wire N__1539;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1524;
    wire N__1521;
    wire N__1518;
    wire N__1515;
    wire N__1512;
    wire N__1509;
    wire N__1506;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1494;
    wire N__1491;
    wire N__1488;
    wire N__1485;
    wire N__1482;
    wire N__1479;
    wire N__1476;
    wire N__1473;
    wire N__1470;
    wire N__1467;
    wire N__1464;
    wire N__1461;
    wire N__1458;
    wire N__1455;
    wire N__1452;
    wire N__1449;
    wire N__1446;
    wire N__1443;
    wire N__1440;
    wire N__1437;
    wire N__1434;
    wire N__1431;
    wire N__1428;
    wire N__1425;
    wire N__1422;
    wire N__1419;
    wire N__1416;
    wire N__1413;
    wire N__1412;
    wire N__1411;
    wire N__1410;
    wire N__1409;
    wire N__1398;
    wire N__1395;
    wire N__1392;
    wire N__1389;
    wire CLK_c_g;
    wire GNDG0;
    wire VCCG0;
    wire CONSTANT_ONE_NET;
    wire SYNTHESIZED_WIRE_4_1;
    wire \b2v_inst3.result_reg1_bmZ0Z_0 ;
    wire \b2v_inst3.result_reg1_amZ0Z_0_cascade_ ;
    wire SYNTHESIZED_WIRE_3_0_cascade_;
    wire N_21;
    wire SYNTHESIZED_WIRE_4_0;
    wire \b2v_inst.A_equal_B_NEZ0Z_2_cascade_ ;
    wire \b2v_inst.A_equal_B_NEZ0Z_0 ;
    wire A_equal_B_c;
    wire SYNTHESIZED_WIRE_0_4_cascade_;
    wire \b2v_inst4.result_reg2_bmZ0Z_4_cascade_ ;
    wire SYNTHESIZED_WIRE_4_4;
    wire SYNTHESIZED_WIRE_0_5_cascade_;
    wire \b2v_inst4.result_reg2_bmZ0Z_5_cascade_ ;
    wire SYNTHESIZED_WIRE_4_5;
    wire N_22;
    wire N_24_cascade_;
    wire SYNTHESIZED_WIRE_4_3;
    wire \b2v_inst4.result_reg2_amZ0Z_4 ;
    wire \b2v_inst4.result_reg2_amZ0Z_5 ;
    wire \b2v_inst4.result_reg2_amZ0Z_7_cascade_ ;
    wire SYNTHESIZED_WIRE_4_7;
    wire bfn_1_11_0_;
    wire \b2v_inst.result_arith_1_1 ;
    wire \b2v_inst.result_arith_1_cry_0 ;
    wire \b2v_inst.result_arith_1_cry_1 ;
    wire \b2v_inst.result_arith_1_3 ;
    wire \b2v_inst.result_arith_1_cry_2 ;
    wire b2v_inst_result_arith_1_4;
    wire \b2v_inst.result_arith_1_cry_3 ;
    wire b2v_inst_result_arith_1_5;
    wire \b2v_inst.result_arith_1_cry_4 ;
    wire \b2v_inst.result_arith_1_cry_5 ;
    wire b2v_inst_result_arith_1_7;
    wire \b2v_inst.result_arith_1_cry_6 ;
    wire \b2v_inst.result_arith_1_8 ;
    wire bfn_1_12_0_;
    wire carry_out_c;
    wire \b2v_inst.A_c_i_0 ;
    wire bfn_1_13_0_;
    wire \b2v_inst.A_c_i_1 ;
    wire \b2v_inst.B_bigger_cry_0 ;
    wire \b2v_inst.A_c_i_2 ;
    wire \b2v_inst.B_bigger_cry_1 ;
    wire \b2v_inst.A_c_i_3 ;
    wire \b2v_inst.B_bigger_cry_2 ;
    wire \b2v_inst.A_c_i_4 ;
    wire \b2v_inst.B_bigger_cry_3 ;
    wire \b2v_inst.A_c_i_5 ;
    wire \b2v_inst.B_bigger_cry_4 ;
    wire \b2v_inst.A_c_i_6 ;
    wire \b2v_inst.B_bigger_cry_5 ;
    wire \b2v_inst.A_c_i_7 ;
    wire \b2v_inst.B_bigger_cry_6 ;
    wire B_bigger_c;
    wire bfn_1_14_0_;
    wire B_bigger_c_THRU_CO;
    wire \b2v_inst3.result_reg1_amZ0Z_1_cascade_ ;
    wire \b2v_inst3.result_reg1_bmZ0Z_1 ;
    wire SYNTHESIZED_WIRE_3_1;
    wire \b2v_inst3.result_reg1_bmZ0Z_3_cascade_ ;
    wire SYNTHESIZED_WIRE_3_3;
    wire \b2v_inst3.result_reg1_amZ0Z_3 ;
    wire \b2v_inst.A_equal_B_NEZ0Z_1 ;
    wire \b2v_inst3.result_reg1_bmZ0Z_2_cascade_ ;
    wire \b2v_inst3.result_reg1_amZ0Z_2 ;
    wire SYNTHESIZED_WIRE_3_2_cascade_;
    wire SYNTHESIZED_WIRE_4_2;
    wire \b2v_inst.A_equal_B_NEZ0Z_3 ;
    wire \b2v_inst.result_arith_1_2 ;
    wire N_23;
    wire s2_c;
    wire SYNTHESIZED_WIRE_4_6;
    wire SYNTHESIZED_WIRE_0_7_cascade_;
    wire \b2v_inst4.result_reg2_bmZ0Z_7 ;
    wire b2v_inst_result_arith_1_6;
    wire \b2v_inst4.result_reg2_amZ0Z_6 ;
    wire S2_S3_c_0;
    wire S2_S3_c_1;
    wire SYNTHESIZED_WIRE_0_6_cascade_;
    wire S1_c;
    wire \b2v_inst4.result_reg2_bmZ0Z_6 ;
    wire bfn_2_11_0_;
    wire \b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4 ;
    wire \b2v_inst.un8_result_arith_cry_0 ;
    wire \b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4 ;
    wire \b2v_inst.un8_result_arith_cry_1 ;
    wire \b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4 ;
    wire \b2v_inst.un8_result_arith_cry_2 ;
    wire un8_result_arith_cry_3_c_RNIO6R4;
    wire \b2v_inst.un8_result_arith_cry_3 ;
    wire un8_result_arith_cry_4_c_RNIQ9S4;
    wire \b2v_inst.un8_result_arith_cry_4 ;
    wire un8_result_arith_cry_5_c_RNISCT4;
    wire \b2v_inst.un8_result_arith_cry_5 ;
    wire \b2v_inst.un8_result_arith_cry_6 ;
    wire un8_result_arith_cry_6_c_RNIK5GH;
    wire B_c_0;
    wire A_c_0;
    wire \b2v_inst.B_c_i_0 ;
    wire bfn_2_12_0_;
    wire A_c_1;
    wire B_c_1;
    wire \b2v_inst.B_c_i_1 ;
    wire \b2v_inst.A_bigger_cry_0 ;
    wire A_c_2;
    wire B_c_2;
    wire \b2v_inst.B_c_i_2 ;
    wire \b2v_inst.A_bigger_cry_1 ;
    wire B_c_3;
    wire A_c_3;
    wire \b2v_inst.B_c_i_3 ;
    wire \b2v_inst.A_bigger_cry_2 ;
    wire A_c_4;
    wire B_c_4;
    wire \b2v_inst.B_c_i_4 ;
    wire \b2v_inst.A_bigger_cry_3 ;
    wire B_c_5;
    wire A_c_5;
    wire \b2v_inst.B_c_i_5 ;
    wire \b2v_inst.A_bigger_cry_4 ;
    wire B_c_6;
    wire A_c_6;
    wire \b2v_inst.B_c_i_6 ;
    wire \b2v_inst.A_bigger_cry_5 ;
    wire B_c_7;
    wire A_c_7;
    wire \b2v_inst.B_c_i_7 ;
    wire \b2v_inst.A_bigger_cry_6 ;
    wire A_bigger_c;
    wire bfn_2_13_0_;
    wire A_bigger_c_THRU_CO;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3706),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__3708),
            .DIN(N__3707),
            .DOUT(N__3706),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__3708),
            .PADOUT(N__3707),
            .PADIN(N__3706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__3697),
            .DIN(N__3696),
            .DOUT(N__3695),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__3697),
            .PADOUT(N__3696),
            .PADIN(N__3695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_7_iopad (
            .OE(N__3688),
            .DIN(N__3687),
            .DOUT(N__3686),
            .PACKAGEPIN(B[7]));
    defparam B_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_7_preio (
            .PADOEN(N__3688),
            .PADOUT(N__3687),
            .PADIN(N__3686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__3679),
            .DIN(N__3678),
            .DOUT(N__3677),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__3679),
            .PADOUT(N__3678),
            .PADIN(N__3677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_6_iopad (
            .OE(N__3670),
            .DIN(N__3669),
            .DOUT(N__3668),
            .PACKAGEPIN(B[6]));
    defparam B_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_6_preio (
            .PADOEN(N__3670),
            .PADOUT(N__3669),
            .PADIN(N__3668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_2_iopad (
            .OE(N__3661),
            .DIN(N__3660),
            .DOUT(N__3659),
            .PACKAGEPIN(F[2]));
    defparam F_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_2_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_2_preio (
            .PADOEN(N__3661),
            .PADOUT(N__3660),
            .PADIN(N__3659),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1412));
    IO_PAD A_ibuf_7_iopad (
            .OE(N__3652),
            .DIN(N__3651),
            .DOUT(N__3650),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__3652),
            .PADOUT(N__3651),
            .PADIN(N__3650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_2_iopad (
            .OE(N__3643),
            .DIN(N__3642),
            .DOUT(N__3641),
            .PACKAGEPIN(B[2]));
    defparam B_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_2_preio (
            .PADOEN(N__3643),
            .PADOUT(N__3642),
            .PADIN(N__3641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_5_iopad (
            .OE(N__3634),
            .DIN(N__3633),
            .DOUT(N__3632),
            .PACKAGEPIN(F[5]));
    defparam F_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_5_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_5_preio (
            .PADOEN(N__3634),
            .PADOUT(N__3633),
            .PADIN(N__3632),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1530),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1409));
    IO_PAD S2_S3_ibuf_0_iopad (
            .OE(N__3625),
            .DIN(N__3624),
            .DOUT(N__3623),
            .PACKAGEPIN(S2_S3[0]));
    defparam S2_S3_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam S2_S3_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO S2_S3_ibuf_0_preio (
            .PADOEN(N__3625),
            .PADOUT(N__3624),
            .PADIN(N__3623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(S2_S3_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD carry_out_obuf_iopad (
            .OE(N__3616),
            .DIN(N__3615),
            .DOUT(N__3614),
            .PACKAGEPIN(carry_out));
    defparam carry_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam carry_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO carry_out_obuf_preio (
            .PADOEN(N__3616),
            .PADOUT(N__3615),
            .PADIN(N__3614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD flag_zero_obuf_iopad (
            .OE(N__3607),
            .DIN(N__3606),
            .DOUT(N__3605),
            .PACKAGEPIN(flag_zero));
    defparam flag_zero_obuf_preio.NEG_TRIGGER=1'b0;
    defparam flag_zero_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO flag_zero_obuf_preio (
            .PADOEN(N__3607),
            .PADOUT(N__3606),
            .PADIN(N__3605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1392),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_1_iopad (
            .OE(N__3598),
            .DIN(N__3597),
            .DOUT(N__3596),
            .PACKAGEPIN(F[1]));
    defparam F_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_1_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_1_preio (
            .PADOEN(N__3598),
            .PADOUT(N__3597),
            .PADIN(N__3596),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1413));
    IO_PAD A_ibuf_0_iopad (
            .OE(N__3589),
            .DIN(N__3588),
            .DOUT(N__3587),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__3589),
            .PADOUT(N__3588),
            .PADIN(N__3587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_5_iopad (
            .OE(N__3580),
            .DIN(N__3579),
            .DOUT(N__3578),
            .PACKAGEPIN(B[5]));
    defparam B_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_5_preio (
            .PADOEN(N__3580),
            .PADOUT(N__3579),
            .PADIN(N__3578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_4_iopad (
            .OE(N__3571),
            .DIN(N__3570),
            .DOUT(N__3569),
            .PACKAGEPIN(F[4]));
    defparam F_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_4_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_4_preio (
            .PADOEN(N__3571),
            .PADOUT(N__3570),
            .PADIN(N__3569),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1411));
    IO_PAD A_equal_B_obuf_iopad (
            .OE(N__3562),
            .DIN(N__3561),
            .DOUT(N__3560),
            .PACKAGEPIN(A_equal_B));
    defparam A_equal_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A_equal_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A_equal_B_obuf_preio (
            .PADOEN(N__3562),
            .PADOUT(N__3561),
            .PADIN(N__3560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD S1_ibuf_iopad (
            .OE(N__3553),
            .DIN(N__3552),
            .DOUT(N__3551),
            .PACKAGEPIN(S1));
    defparam S1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam S1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO S1_ibuf_preio (
            .PADOEN(N__3553),
            .PADOUT(N__3552),
            .PADIN(N__3551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(S1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__3544),
            .DIN(N__3543),
            .DOUT(N__3542),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__3544),
            .PADOUT(N__3543),
            .PADIN(N__3542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_1_iopad (
            .OE(N__3535),
            .DIN(N__3534),
            .DOUT(N__3533),
            .PACKAGEPIN(B[1]));
    defparam B_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_1_preio (
            .PADOEN(N__3535),
            .PADOUT(N__3534),
            .PADIN(N__3533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_0_iopad (
            .OE(N__3526),
            .DIN(N__3525),
            .DOUT(N__3524),
            .PACKAGEPIN(F[0]));
    defparam F_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_0_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_0_preio (
            .PADOEN(N__3526),
            .PADOUT(N__3525),
            .PADIN(N__3524),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1411));
    IO_PAD s2_ibuf_iopad (
            .OE(N__3517),
            .DIN(N__3516),
            .DOUT(N__3515),
            .PACKAGEPIN(s2));
    defparam s2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO s2_ibuf_preio (
            .PADOEN(N__3517),
            .PADOUT(N__3516),
            .PADIN(N__3515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(s2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_bigger_obuf_iopad (
            .OE(N__3508),
            .DIN(N__3507),
            .DOUT(N__3506),
            .PACKAGEPIN(B_bigger));
    defparam B_bigger_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_bigger_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_bigger_obuf_preio (
            .PADOEN(N__3508),
            .PADOUT(N__3507),
            .PADIN(N__3506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1731),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__3499),
            .DIN(N__3498),
            .DOUT(N__3497),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__3499),
            .PADOUT(N__3498),
            .PADIN(N__3497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_4_iopad (
            .OE(N__3490),
            .DIN(N__3489),
            .DOUT(N__3488),
            .PACKAGEPIN(B[4]));
    defparam B_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_4_preio (
            .PADOEN(N__3490),
            .PADOUT(N__3489),
            .PADIN(N__3488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD over_flow_obuf_iopad (
            .OE(N__3481),
            .DIN(N__3480),
            .DOUT(N__3479),
            .PACKAGEPIN(over_flow));
    defparam over_flow_obuf_preio.NEG_TRIGGER=1'b0;
    defparam over_flow_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO over_flow_obuf_preio (
            .PADOEN(N__3481),
            .PADOUT(N__3480),
            .PADIN(N__3479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__3472),
            .DIN(N__3471),
            .DOUT(N__3470),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__3472),
            .PADOUT(N__3471),
            .PADIN(N__3470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_0_iopad (
            .OE(N__3463),
            .DIN(N__3462),
            .DOUT(N__3461),
            .PACKAGEPIN(B[0]));
    defparam B_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_0_preio (
            .PADOEN(N__3463),
            .PADOUT(N__3462),
            .PADIN(N__3461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_7_iopad (
            .OE(N__3454),
            .DIN(N__3453),
            .DOUT(N__3452),
            .PACKAGEPIN(F[7]));
    defparam F_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_7_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_7_preio (
            .PADOEN(N__3454),
            .PADOUT(N__3453),
            .PADIN(N__3452),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1605),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1410));
    IO_PAD A_bigger_obuf_iopad (
            .OE(N__3445),
            .DIN(N__3444),
            .DOUT(N__3443),
            .PACKAGEPIN(A_bigger));
    defparam A_bigger_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A_bigger_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A_bigger_obuf_preio (
            .PADOEN(N__3445),
            .PADOUT(N__3444),
            .PADIN(N__3443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_3_iopad (
            .OE(N__3436),
            .DIN(N__3435),
            .DOUT(N__3434),
            .PACKAGEPIN(F[3]));
    defparam F_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_3_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_3_preio (
            .PADOEN(N__3436),
            .PADOUT(N__3435),
            .PADIN(N__3434),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1509),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1412));
    IO_PAD A_ibuf_6_iopad (
            .OE(N__3427),
            .DIN(N__3426),
            .DOUT(N__3425),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__3427),
            .PADOUT(N__3426),
            .PADIN(N__3425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_3_iopad (
            .OE(N__3418),
            .DIN(N__3417),
            .DOUT(N__3416),
            .PACKAGEPIN(B[3]));
    defparam B_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_3_preio (
            .PADOEN(N__3418),
            .PADOUT(N__3417),
            .PADIN(N__3416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_obuf_6_iopad (
            .OE(N__3409),
            .DIN(N__3408),
            .DOUT(N__3407),
            .PACKAGEPIN(F[6]));
    defparam F_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam F_obuf_6_preio.PIN_TYPE=6'b010101;
    PRE_IO F_obuf_6_preio (
            .PADOEN(N__3409),
            .PADOUT(N__3408),
            .PADIN(N__3407),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1755),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1410));
    IO_PAD S2_S3_ibuf_1_iopad (
            .OE(N__3400),
            .DIN(N__3399),
            .DOUT(N__3398),
            .PACKAGEPIN(S2_S3[1]));
    defparam S2_S3_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam S2_S3_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO S2_S3_ibuf_1_preio (
            .PADOEN(N__3400),
            .PADOUT(N__3399),
            .PADIN(N__3398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(S2_S3_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__786 (
            .O(N__3381),
            .I(N__3370));
    InMux I__785 (
            .O(N__3380),
            .I(N__3370));
    InMux I__784 (
            .O(N__3379),
            .I(N__3370));
    CascadeMux I__783 (
            .O(N__3378),
            .I(N__3366));
    CascadeMux I__782 (
            .O(N__3377),
            .I(N__3363));
    LocalMux I__781 (
            .O(N__3370),
            .I(N__3360));
    InMux I__780 (
            .O(N__3369),
            .I(N__3357));
    InMux I__779 (
            .O(N__3366),
            .I(N__3354));
    InMux I__778 (
            .O(N__3363),
            .I(N__3351));
    Span4Mux_s1_h I__777 (
            .O(N__3360),
            .I(N__3344));
    LocalMux I__776 (
            .O(N__3357),
            .I(N__3344));
    LocalMux I__775 (
            .O(N__3354),
            .I(N__3344));
    LocalMux I__774 (
            .O(N__3351),
            .I(N__3341));
    Span4Mux_v I__773 (
            .O(N__3344),
            .I(N__3337));
    Span4Mux_v I__772 (
            .O(N__3341),
            .I(N__3334));
    InMux I__771 (
            .O(N__3340),
            .I(N__3331));
    Odrv4 I__770 (
            .O(N__3337),
            .I(A_c_4));
    Odrv4 I__769 (
            .O(N__3334),
            .I(A_c_4));
    LocalMux I__768 (
            .O(N__3331),
            .I(A_c_4));
    CascadeMux I__767 (
            .O(N__3324),
            .I(N__3319));
    CascadeMux I__766 (
            .O(N__3323),
            .I(N__3316));
    InMux I__765 (
            .O(N__3322),
            .I(N__3311));
    InMux I__764 (
            .O(N__3319),
            .I(N__3311));
    InMux I__763 (
            .O(N__3316),
            .I(N__3308));
    LocalMux I__762 (
            .O(N__3311),
            .I(N__3303));
    LocalMux I__761 (
            .O(N__3308),
            .I(N__3300));
    InMux I__760 (
            .O(N__3307),
            .I(N__3297));
    InMux I__759 (
            .O(N__3306),
            .I(N__3294));
    Span4Mux_v I__758 (
            .O(N__3303),
            .I(N__3289));
    Span4Mux_v I__757 (
            .O(N__3300),
            .I(N__3289));
    LocalMux I__756 (
            .O(N__3297),
            .I(N__3286));
    LocalMux I__755 (
            .O(N__3294),
            .I(B_c_4));
    Odrv4 I__754 (
            .O(N__3289),
            .I(B_c_4));
    Odrv4 I__753 (
            .O(N__3286),
            .I(B_c_4));
    CascadeMux I__752 (
            .O(N__3279),
            .I(N__3276));
    InMux I__751 (
            .O(N__3276),
            .I(N__3272));
    InMux I__750 (
            .O(N__3275),
            .I(N__3269));
    LocalMux I__749 (
            .O(N__3272),
            .I(\b2v_inst.B_c_i_4 ));
    LocalMux I__748 (
            .O(N__3269),
            .I(\b2v_inst.B_c_i_4 ));
    InMux I__747 (
            .O(N__3264),
            .I(N__3258));
    InMux I__746 (
            .O(N__3263),
            .I(N__3258));
    LocalMux I__745 (
            .O(N__3258),
            .I(N__3253));
    CascadeMux I__744 (
            .O(N__3257),
            .I(N__3249));
    InMux I__743 (
            .O(N__3256),
            .I(N__3246));
    Span4Mux_v I__742 (
            .O(N__3253),
            .I(N__3243));
    InMux I__741 (
            .O(N__3252),
            .I(N__3240));
    InMux I__740 (
            .O(N__3249),
            .I(N__3237));
    LocalMux I__739 (
            .O(N__3246),
            .I(N__3234));
    Odrv4 I__738 (
            .O(N__3243),
            .I(B_c_5));
    LocalMux I__737 (
            .O(N__3240),
            .I(B_c_5));
    LocalMux I__736 (
            .O(N__3237),
            .I(B_c_5));
    Odrv12 I__735 (
            .O(N__3234),
            .I(B_c_5));
    CascadeMux I__734 (
            .O(N__3225),
            .I(N__3218));
    CascadeMux I__733 (
            .O(N__3224),
            .I(N__3214));
    InMux I__732 (
            .O(N__3223),
            .I(N__3211));
    CascadeMux I__731 (
            .O(N__3222),
            .I(N__3208));
    CascadeMux I__730 (
            .O(N__3221),
            .I(N__3205));
    InMux I__729 (
            .O(N__3218),
            .I(N__3200));
    InMux I__728 (
            .O(N__3217),
            .I(N__3200));
    InMux I__727 (
            .O(N__3214),
            .I(N__3196));
    LocalMux I__726 (
            .O(N__3211),
            .I(N__3193));
    InMux I__725 (
            .O(N__3208),
            .I(N__3190));
    InMux I__724 (
            .O(N__3205),
            .I(N__3187));
    LocalMux I__723 (
            .O(N__3200),
            .I(N__3184));
    InMux I__722 (
            .O(N__3199),
            .I(N__3181));
    LocalMux I__721 (
            .O(N__3196),
            .I(N__3178));
    Span4Mux_s3_h I__720 (
            .O(N__3193),
            .I(N__3175));
    LocalMux I__719 (
            .O(N__3190),
            .I(N__3170));
    LocalMux I__718 (
            .O(N__3187),
            .I(N__3170));
    Span4Mux_s3_h I__717 (
            .O(N__3184),
            .I(N__3167));
    LocalMux I__716 (
            .O(N__3181),
            .I(N__3164));
    Span4Mux_s3_h I__715 (
            .O(N__3178),
            .I(N__3161));
    Span4Mux_v I__714 (
            .O(N__3175),
            .I(N__3158));
    Span12Mux_s3_h I__713 (
            .O(N__3170),
            .I(N__3155));
    Span4Mux_v I__712 (
            .O(N__3167),
            .I(N__3150));
    Span4Mux_s3_h I__711 (
            .O(N__3164),
            .I(N__3150));
    Span4Mux_v I__710 (
            .O(N__3161),
            .I(N__3147));
    Odrv4 I__709 (
            .O(N__3158),
            .I(A_c_5));
    Odrv12 I__708 (
            .O(N__3155),
            .I(A_c_5));
    Odrv4 I__707 (
            .O(N__3150),
            .I(A_c_5));
    Odrv4 I__706 (
            .O(N__3147),
            .I(A_c_5));
    InMux I__705 (
            .O(N__3138),
            .I(N__3134));
    InMux I__704 (
            .O(N__3137),
            .I(N__3131));
    LocalMux I__703 (
            .O(N__3134),
            .I(\b2v_inst.B_c_i_5 ));
    LocalMux I__702 (
            .O(N__3131),
            .I(\b2v_inst.B_c_i_5 ));
    InMux I__701 (
            .O(N__3126),
            .I(N__3118));
    InMux I__700 (
            .O(N__3125),
            .I(N__3118));
    InMux I__699 (
            .O(N__3124),
            .I(N__3115));
    InMux I__698 (
            .O(N__3123),
            .I(N__3112));
    LocalMux I__697 (
            .O(N__3118),
            .I(N__3104));
    LocalMux I__696 (
            .O(N__3115),
            .I(N__3104));
    LocalMux I__695 (
            .O(N__3112),
            .I(N__3104));
    CascadeMux I__694 (
            .O(N__3111),
            .I(N__3101));
    Span4Mux_v I__693 (
            .O(N__3104),
            .I(N__3098));
    InMux I__692 (
            .O(N__3101),
            .I(N__3095));
    Odrv4 I__691 (
            .O(N__3098),
            .I(B_c_6));
    LocalMux I__690 (
            .O(N__3095),
            .I(B_c_6));
    CascadeMux I__689 (
            .O(N__3090),
            .I(N__3085));
    InMux I__688 (
            .O(N__3089),
            .I(N__3075));
    InMux I__687 (
            .O(N__3088),
            .I(N__3075));
    InMux I__686 (
            .O(N__3085),
            .I(N__3075));
    CascadeMux I__685 (
            .O(N__3084),
            .I(N__3072));
    CascadeMux I__684 (
            .O(N__3083),
            .I(N__3069));
    CascadeMux I__683 (
            .O(N__3082),
            .I(N__3066));
    LocalMux I__682 (
            .O(N__3075),
            .I(N__3063));
    InMux I__681 (
            .O(N__3072),
            .I(N__3060));
    InMux I__680 (
            .O(N__3069),
            .I(N__3057));
    InMux I__679 (
            .O(N__3066),
            .I(N__3054));
    Span4Mux_h I__678 (
            .O(N__3063),
            .I(N__3047));
    LocalMux I__677 (
            .O(N__3060),
            .I(N__3047));
    LocalMux I__676 (
            .O(N__3057),
            .I(N__3047));
    LocalMux I__675 (
            .O(N__3054),
            .I(N__3044));
    Span4Mux_v I__674 (
            .O(N__3047),
            .I(N__3040));
    Span4Mux_v I__673 (
            .O(N__3044),
            .I(N__3037));
    InMux I__672 (
            .O(N__3043),
            .I(N__3034));
    Odrv4 I__671 (
            .O(N__3040),
            .I(A_c_6));
    Odrv4 I__670 (
            .O(N__3037),
            .I(A_c_6));
    LocalMux I__669 (
            .O(N__3034),
            .I(A_c_6));
    InMux I__668 (
            .O(N__3027),
            .I(N__3023));
    InMux I__667 (
            .O(N__3026),
            .I(N__3020));
    LocalMux I__666 (
            .O(N__3023),
            .I(\b2v_inst.B_c_i_6 ));
    LocalMux I__665 (
            .O(N__3020),
            .I(\b2v_inst.B_c_i_6 ));
    InMux I__664 (
            .O(N__3015),
            .I(N__3007));
    InMux I__663 (
            .O(N__3014),
            .I(N__3007));
    InMux I__662 (
            .O(N__3013),
            .I(N__3004));
    InMux I__661 (
            .O(N__3012),
            .I(N__3001));
    LocalMux I__660 (
            .O(N__3007),
            .I(N__2997));
    LocalMux I__659 (
            .O(N__3004),
            .I(N__2994));
    LocalMux I__658 (
            .O(N__3001),
            .I(N__2991));
    CascadeMux I__657 (
            .O(N__3000),
            .I(N__2987));
    Span4Mux_h I__656 (
            .O(N__2997),
            .I(N__2984));
    Span4Mux_h I__655 (
            .O(N__2994),
            .I(N__2981));
    Span4Mux_h I__654 (
            .O(N__2991),
            .I(N__2978));
    InMux I__653 (
            .O(N__2990),
            .I(N__2975));
    InMux I__652 (
            .O(N__2987),
            .I(N__2972));
    Span4Mux_v I__651 (
            .O(N__2984),
            .I(N__2969));
    Span4Mux_v I__650 (
            .O(N__2981),
            .I(N__2966));
    Sp12to4 I__649 (
            .O(N__2978),
            .I(N__2959));
    LocalMux I__648 (
            .O(N__2975),
            .I(N__2959));
    LocalMux I__647 (
            .O(N__2972),
            .I(N__2959));
    Odrv4 I__646 (
            .O(N__2969),
            .I(B_c_7));
    Odrv4 I__645 (
            .O(N__2966),
            .I(B_c_7));
    Odrv12 I__644 (
            .O(N__2959),
            .I(B_c_7));
    CascadeMux I__643 (
            .O(N__2952),
            .I(N__2949));
    InMux I__642 (
            .O(N__2949),
            .I(N__2941));
    InMux I__641 (
            .O(N__2948),
            .I(N__2941));
    CascadeMux I__640 (
            .O(N__2947),
            .I(N__2938));
    CascadeMux I__639 (
            .O(N__2946),
            .I(N__2934));
    LocalMux I__638 (
            .O(N__2941),
            .I(N__2931));
    InMux I__637 (
            .O(N__2938),
            .I(N__2928));
    InMux I__636 (
            .O(N__2937),
            .I(N__2925));
    InMux I__635 (
            .O(N__2934),
            .I(N__2922));
    Span4Mux_h I__634 (
            .O(N__2931),
            .I(N__2917));
    LocalMux I__633 (
            .O(N__2928),
            .I(N__2917));
    LocalMux I__632 (
            .O(N__2925),
            .I(N__2914));
    LocalMux I__631 (
            .O(N__2922),
            .I(N__2911));
    Span4Mux_v I__630 (
            .O(N__2917),
            .I(N__2907));
    Span4Mux_v I__629 (
            .O(N__2914),
            .I(N__2902));
    Span4Mux_v I__628 (
            .O(N__2911),
            .I(N__2902));
    InMux I__627 (
            .O(N__2910),
            .I(N__2899));
    Odrv4 I__626 (
            .O(N__2907),
            .I(A_c_7));
    Odrv4 I__625 (
            .O(N__2902),
            .I(A_c_7));
    LocalMux I__624 (
            .O(N__2899),
            .I(A_c_7));
    InMux I__623 (
            .O(N__2892),
            .I(N__2889));
    LocalMux I__622 (
            .O(N__2889),
            .I(\b2v_inst.B_c_i_7 ));
    InMux I__621 (
            .O(N__2886),
            .I(bfn_2_13_0_));
    IoInMux I__620 (
            .O(N__2883),
            .I(N__2880));
    LocalMux I__619 (
            .O(N__2880),
            .I(N__2877));
    Span4Mux_s3_v I__618 (
            .O(N__2877),
            .I(N__2874));
    Odrv4 I__617 (
            .O(N__2874),
            .I(A_bigger_c_THRU_CO));
    InMux I__616 (
            .O(N__2871),
            .I(N__2868));
    LocalMux I__615 (
            .O(N__2868),
            .I(un8_result_arith_cry_4_c_RNIQ9S4));
    InMux I__614 (
            .O(N__2865),
            .I(\b2v_inst.un8_result_arith_cry_4 ));
    InMux I__613 (
            .O(N__2862),
            .I(N__2859));
    LocalMux I__612 (
            .O(N__2859),
            .I(un8_result_arith_cry_5_c_RNISCT4));
    InMux I__611 (
            .O(N__2856),
            .I(\b2v_inst.un8_result_arith_cry_5 ));
    InMux I__610 (
            .O(N__2853),
            .I(\b2v_inst.un8_result_arith_cry_6 ));
    InMux I__609 (
            .O(N__2850),
            .I(N__2847));
    LocalMux I__608 (
            .O(N__2847),
            .I(un8_result_arith_cry_6_c_RNIK5GH));
    CascadeMux I__607 (
            .O(N__2844),
            .I(N__2839));
    CascadeMux I__606 (
            .O(N__2843),
            .I(N__2835));
    CascadeMux I__605 (
            .O(N__2842),
            .I(N__2832));
    InMux I__604 (
            .O(N__2839),
            .I(N__2828));
    InMux I__603 (
            .O(N__2838),
            .I(N__2823));
    InMux I__602 (
            .O(N__2835),
            .I(N__2823));
    InMux I__601 (
            .O(N__2832),
            .I(N__2820));
    InMux I__600 (
            .O(N__2831),
            .I(N__2817));
    LocalMux I__599 (
            .O(N__2828),
            .I(N__2814));
    LocalMux I__598 (
            .O(N__2823),
            .I(N__2811));
    LocalMux I__597 (
            .O(N__2820),
            .I(N__2806));
    LocalMux I__596 (
            .O(N__2817),
            .I(N__2806));
    Span4Mux_v I__595 (
            .O(N__2814),
            .I(N__2798));
    Span4Mux_v I__594 (
            .O(N__2811),
            .I(N__2798));
    Span4Mux_v I__593 (
            .O(N__2806),
            .I(N__2798));
    InMux I__592 (
            .O(N__2805),
            .I(N__2795));
    Odrv4 I__591 (
            .O(N__2798),
            .I(B_c_0));
    LocalMux I__590 (
            .O(N__2795),
            .I(B_c_0));
    CascadeMux I__589 (
            .O(N__2790),
            .I(N__2787));
    InMux I__588 (
            .O(N__2787),
            .I(N__2775));
    InMux I__587 (
            .O(N__2786),
            .I(N__2775));
    InMux I__586 (
            .O(N__2785),
            .I(N__2775));
    InMux I__585 (
            .O(N__2784),
            .I(N__2772));
    CascadeMux I__584 (
            .O(N__2783),
            .I(N__2767));
    CascadeMux I__583 (
            .O(N__2782),
            .I(N__2764));
    LocalMux I__582 (
            .O(N__2775),
            .I(N__2761));
    LocalMux I__581 (
            .O(N__2772),
            .I(N__2758));
    InMux I__580 (
            .O(N__2771),
            .I(N__2755));
    CascadeMux I__579 (
            .O(N__2770),
            .I(N__2752));
    InMux I__578 (
            .O(N__2767),
            .I(N__2748));
    InMux I__577 (
            .O(N__2764),
            .I(N__2745));
    Span4Mux_s2_h I__576 (
            .O(N__2761),
            .I(N__2741));
    Span4Mux_s2_h I__575 (
            .O(N__2758),
            .I(N__2738));
    LocalMux I__574 (
            .O(N__2755),
            .I(N__2735));
    InMux I__573 (
            .O(N__2752),
            .I(N__2732));
    InMux I__572 (
            .O(N__2751),
            .I(N__2729));
    LocalMux I__571 (
            .O(N__2748),
            .I(N__2726));
    LocalMux I__570 (
            .O(N__2745),
            .I(N__2723));
    InMux I__569 (
            .O(N__2744),
            .I(N__2720));
    Span4Mux_v I__568 (
            .O(N__2741),
            .I(N__2715));
    Span4Mux_v I__567 (
            .O(N__2738),
            .I(N__2715));
    Span4Mux_v I__566 (
            .O(N__2735),
            .I(N__2710));
    LocalMux I__565 (
            .O(N__2732),
            .I(N__2710));
    LocalMux I__564 (
            .O(N__2729),
            .I(N__2707));
    Span4Mux_v I__563 (
            .O(N__2726),
            .I(N__2700));
    Span4Mux_s2_h I__562 (
            .O(N__2723),
            .I(N__2700));
    LocalMux I__561 (
            .O(N__2720),
            .I(N__2700));
    Span4Mux_v I__560 (
            .O(N__2715),
            .I(N__2697));
    Span4Mux_v I__559 (
            .O(N__2710),
            .I(N__2692));
    Span4Mux_s2_h I__558 (
            .O(N__2707),
            .I(N__2692));
    Span4Mux_v I__557 (
            .O(N__2700),
            .I(N__2689));
    Odrv4 I__556 (
            .O(N__2697),
            .I(A_c_0));
    Odrv4 I__555 (
            .O(N__2692),
            .I(A_c_0));
    Odrv4 I__554 (
            .O(N__2689),
            .I(A_c_0));
    CascadeMux I__553 (
            .O(N__2682),
            .I(N__2678));
    InMux I__552 (
            .O(N__2681),
            .I(N__2675));
    InMux I__551 (
            .O(N__2678),
            .I(N__2672));
    LocalMux I__550 (
            .O(N__2675),
            .I(\b2v_inst.B_c_i_0 ));
    LocalMux I__549 (
            .O(N__2672),
            .I(\b2v_inst.B_c_i_0 ));
    InMux I__548 (
            .O(N__2667),
            .I(N__2658));
    InMux I__547 (
            .O(N__2666),
            .I(N__2658));
    CascadeMux I__546 (
            .O(N__2665),
            .I(N__2654));
    CascadeMux I__545 (
            .O(N__2664),
            .I(N__2651));
    CascadeMux I__544 (
            .O(N__2663),
            .I(N__2647));
    LocalMux I__543 (
            .O(N__2658),
            .I(N__2644));
    InMux I__542 (
            .O(N__2657),
            .I(N__2640));
    InMux I__541 (
            .O(N__2654),
            .I(N__2637));
    InMux I__540 (
            .O(N__2651),
            .I(N__2634));
    CascadeMux I__539 (
            .O(N__2650),
            .I(N__2631));
    InMux I__538 (
            .O(N__2647),
            .I(N__2628));
    Span4Mux_v I__537 (
            .O(N__2644),
            .I(N__2625));
    InMux I__536 (
            .O(N__2643),
            .I(N__2622));
    LocalMux I__535 (
            .O(N__2640),
            .I(N__2617));
    LocalMux I__534 (
            .O(N__2637),
            .I(N__2617));
    LocalMux I__533 (
            .O(N__2634),
            .I(N__2614));
    InMux I__532 (
            .O(N__2631),
            .I(N__2611));
    LocalMux I__531 (
            .O(N__2628),
            .I(N__2608));
    Span4Mux_v I__530 (
            .O(N__2625),
            .I(N__2605));
    LocalMux I__529 (
            .O(N__2622),
            .I(N__2602));
    Span4Mux_v I__528 (
            .O(N__2617),
            .I(N__2595));
    Span4Mux_s2_h I__527 (
            .O(N__2614),
            .I(N__2595));
    LocalMux I__526 (
            .O(N__2611),
            .I(N__2595));
    Span4Mux_v I__525 (
            .O(N__2608),
            .I(N__2592));
    IoSpan4Mux I__524 (
            .O(N__2605),
            .I(N__2587));
    IoSpan4Mux I__523 (
            .O(N__2602),
            .I(N__2587));
    Span4Mux_v I__522 (
            .O(N__2595),
            .I(N__2584));
    Odrv4 I__521 (
            .O(N__2592),
            .I(A_c_1));
    Odrv4 I__520 (
            .O(N__2587),
            .I(A_c_1));
    Odrv4 I__519 (
            .O(N__2584),
            .I(A_c_1));
    InMux I__518 (
            .O(N__2577),
            .I(N__2571));
    InMux I__517 (
            .O(N__2576),
            .I(N__2568));
    InMux I__516 (
            .O(N__2575),
            .I(N__2565));
    InMux I__515 (
            .O(N__2574),
            .I(N__2562));
    LocalMux I__514 (
            .O(N__2571),
            .I(N__2559));
    LocalMux I__513 (
            .O(N__2568),
            .I(N__2556));
    LocalMux I__512 (
            .O(N__2565),
            .I(N__2553));
    LocalMux I__511 (
            .O(N__2562),
            .I(N__2550));
    Span4Mux_v I__510 (
            .O(N__2559),
            .I(N__2544));
    Span4Mux_v I__509 (
            .O(N__2556),
            .I(N__2544));
    Span4Mux_v I__508 (
            .O(N__2553),
            .I(N__2539));
    Span4Mux_v I__507 (
            .O(N__2550),
            .I(N__2539));
    InMux I__506 (
            .O(N__2549),
            .I(N__2536));
    Odrv4 I__505 (
            .O(N__2544),
            .I(B_c_1));
    Odrv4 I__504 (
            .O(N__2539),
            .I(B_c_1));
    LocalMux I__503 (
            .O(N__2536),
            .I(B_c_1));
    InMux I__502 (
            .O(N__2529),
            .I(N__2525));
    InMux I__501 (
            .O(N__2528),
            .I(N__2522));
    LocalMux I__500 (
            .O(N__2525),
            .I(\b2v_inst.B_c_i_1 ));
    LocalMux I__499 (
            .O(N__2522),
            .I(\b2v_inst.B_c_i_1 ));
    CascadeMux I__498 (
            .O(N__2517),
            .I(N__2512));
    CascadeMux I__497 (
            .O(N__2516),
            .I(N__2508));
    InMux I__496 (
            .O(N__2515),
            .I(N__2505));
    InMux I__495 (
            .O(N__2512),
            .I(N__2502));
    CascadeMux I__494 (
            .O(N__2511),
            .I(N__2498));
    InMux I__493 (
            .O(N__2508),
            .I(N__2495));
    LocalMux I__492 (
            .O(N__2505),
            .I(N__2489));
    LocalMux I__491 (
            .O(N__2502),
            .I(N__2486));
    InMux I__490 (
            .O(N__2501),
            .I(N__2483));
    InMux I__489 (
            .O(N__2498),
            .I(N__2480));
    LocalMux I__488 (
            .O(N__2495),
            .I(N__2477));
    InMux I__487 (
            .O(N__2494),
            .I(N__2470));
    InMux I__486 (
            .O(N__2493),
            .I(N__2470));
    InMux I__485 (
            .O(N__2492),
            .I(N__2470));
    Span4Mux_s1_h I__484 (
            .O(N__2489),
            .I(N__2461));
    Span4Mux_v I__483 (
            .O(N__2486),
            .I(N__2461));
    LocalMux I__482 (
            .O(N__2483),
            .I(N__2461));
    LocalMux I__481 (
            .O(N__2480),
            .I(N__2461));
    Sp12to4 I__480 (
            .O(N__2477),
            .I(N__2456));
    LocalMux I__479 (
            .O(N__2470),
            .I(N__2456));
    Span4Mux_v I__478 (
            .O(N__2461),
            .I(N__2453));
    Odrv12 I__477 (
            .O(N__2456),
            .I(A_c_2));
    Odrv4 I__476 (
            .O(N__2453),
            .I(A_c_2));
    CascadeMux I__475 (
            .O(N__2448),
            .I(N__2443));
    CascadeMux I__474 (
            .O(N__2447),
            .I(N__2440));
    InMux I__473 (
            .O(N__2446),
            .I(N__2437));
    InMux I__472 (
            .O(N__2443),
            .I(N__2431));
    InMux I__471 (
            .O(N__2440),
            .I(N__2431));
    LocalMux I__470 (
            .O(N__2437),
            .I(N__2428));
    CascadeMux I__469 (
            .O(N__2436),
            .I(N__2425));
    LocalMux I__468 (
            .O(N__2431),
            .I(N__2422));
    Span4Mux_h I__467 (
            .O(N__2428),
            .I(N__2418));
    InMux I__466 (
            .O(N__2425),
            .I(N__2415));
    Span4Mux_h I__465 (
            .O(N__2422),
            .I(N__2412));
    InMux I__464 (
            .O(N__2421),
            .I(N__2409));
    Span4Mux_v I__463 (
            .O(N__2418),
            .I(N__2406));
    LocalMux I__462 (
            .O(N__2415),
            .I(N__2403));
    Sp12to4 I__461 (
            .O(N__2412),
            .I(N__2398));
    LocalMux I__460 (
            .O(N__2409),
            .I(N__2398));
    Odrv4 I__459 (
            .O(N__2406),
            .I(B_c_2));
    Odrv12 I__458 (
            .O(N__2403),
            .I(B_c_2));
    Odrv12 I__457 (
            .O(N__2398),
            .I(B_c_2));
    InMux I__456 (
            .O(N__2391),
            .I(N__2387));
    InMux I__455 (
            .O(N__2390),
            .I(N__2384));
    LocalMux I__454 (
            .O(N__2387),
            .I(\b2v_inst.B_c_i_2 ));
    LocalMux I__453 (
            .O(N__2384),
            .I(\b2v_inst.B_c_i_2 ));
    InMux I__452 (
            .O(N__2379),
            .I(N__2374));
    CascadeMux I__451 (
            .O(N__2378),
            .I(N__2371));
    CascadeMux I__450 (
            .O(N__2377),
            .I(N__2368));
    LocalMux I__449 (
            .O(N__2374),
            .I(N__2364));
    InMux I__448 (
            .O(N__2371),
            .I(N__2361));
    InMux I__447 (
            .O(N__2368),
            .I(N__2355));
    InMux I__446 (
            .O(N__2367),
            .I(N__2355));
    Span4Mux_v I__445 (
            .O(N__2364),
            .I(N__2350));
    LocalMux I__444 (
            .O(N__2361),
            .I(N__2350));
    InMux I__443 (
            .O(N__2360),
            .I(N__2347));
    LocalMux I__442 (
            .O(N__2355),
            .I(N__2344));
    Span4Mux_v I__441 (
            .O(N__2350),
            .I(N__2341));
    LocalMux I__440 (
            .O(N__2347),
            .I(N__2338));
    Odrv12 I__439 (
            .O(N__2344),
            .I(B_c_3));
    Odrv4 I__438 (
            .O(N__2341),
            .I(B_c_3));
    Odrv12 I__437 (
            .O(N__2338),
            .I(B_c_3));
    CascadeMux I__436 (
            .O(N__2331),
            .I(N__2325));
    InMux I__435 (
            .O(N__2330),
            .I(N__2315));
    InMux I__434 (
            .O(N__2329),
            .I(N__2315));
    InMux I__433 (
            .O(N__2328),
            .I(N__2315));
    InMux I__432 (
            .O(N__2325),
            .I(N__2312));
    InMux I__431 (
            .O(N__2324),
            .I(N__2308));
    CascadeMux I__430 (
            .O(N__2323),
            .I(N__2305));
    InMux I__429 (
            .O(N__2322),
            .I(N__2302));
    LocalMux I__428 (
            .O(N__2315),
            .I(N__2297));
    LocalMux I__427 (
            .O(N__2312),
            .I(N__2297));
    CascadeMux I__426 (
            .O(N__2311),
            .I(N__2294));
    LocalMux I__425 (
            .O(N__2308),
            .I(N__2291));
    InMux I__424 (
            .O(N__2305),
            .I(N__2288));
    LocalMux I__423 (
            .O(N__2302),
            .I(N__2284));
    Span4Mux_v I__422 (
            .O(N__2297),
            .I(N__2281));
    InMux I__421 (
            .O(N__2294),
            .I(N__2278));
    Span4Mux_s2_h I__420 (
            .O(N__2291),
            .I(N__2273));
    LocalMux I__419 (
            .O(N__2288),
            .I(N__2273));
    InMux I__418 (
            .O(N__2287),
            .I(N__2270));
    Span4Mux_s3_h I__417 (
            .O(N__2284),
            .I(N__2267));
    IoSpan4Mux I__416 (
            .O(N__2281),
            .I(N__2262));
    LocalMux I__415 (
            .O(N__2278),
            .I(N__2262));
    Span4Mux_v I__414 (
            .O(N__2273),
            .I(N__2259));
    LocalMux I__413 (
            .O(N__2270),
            .I(N__2256));
    Span4Mux_v I__412 (
            .O(N__2267),
            .I(N__2251));
    Span4Mux_s3_h I__411 (
            .O(N__2262),
            .I(N__2251));
    IoSpan4Mux I__410 (
            .O(N__2259),
            .I(N__2248));
    Span4Mux_s3_h I__409 (
            .O(N__2256),
            .I(N__2245));
    Span4Mux_v I__408 (
            .O(N__2251),
            .I(N__2242));
    Odrv4 I__407 (
            .O(N__2248),
            .I(A_c_3));
    Odrv4 I__406 (
            .O(N__2245),
            .I(A_c_3));
    Odrv4 I__405 (
            .O(N__2242),
            .I(A_c_3));
    InMux I__404 (
            .O(N__2235),
            .I(N__2231));
    InMux I__403 (
            .O(N__2234),
            .I(N__2228));
    LocalMux I__402 (
            .O(N__2231),
            .I(\b2v_inst.B_c_i_3 ));
    LocalMux I__401 (
            .O(N__2228),
            .I(\b2v_inst.B_c_i_3 ));
    CascadeMux I__400 (
            .O(N__2223),
            .I(SYNTHESIZED_WIRE_0_7_cascade_));
    InMux I__399 (
            .O(N__2220),
            .I(N__2217));
    LocalMux I__398 (
            .O(N__2217),
            .I(\b2v_inst4.result_reg2_bmZ0Z_7 ));
    InMux I__397 (
            .O(N__2214),
            .I(N__2211));
    LocalMux I__396 (
            .O(N__2211),
            .I(b2v_inst_result_arith_1_6));
    InMux I__395 (
            .O(N__2208),
            .I(N__2205));
    LocalMux I__394 (
            .O(N__2205),
            .I(\b2v_inst4.result_reg2_amZ0Z_6 ));
    CascadeMux I__393 (
            .O(N__2202),
            .I(N__2198));
    InMux I__392 (
            .O(N__2201),
            .I(N__2180));
    InMux I__391 (
            .O(N__2198),
            .I(N__2180));
    InMux I__390 (
            .O(N__2197),
            .I(N__2175));
    InMux I__389 (
            .O(N__2196),
            .I(N__2175));
    InMux I__388 (
            .O(N__2195),
            .I(N__2166));
    InMux I__387 (
            .O(N__2194),
            .I(N__2166));
    InMux I__386 (
            .O(N__2193),
            .I(N__2166));
    InMux I__385 (
            .O(N__2192),
            .I(N__2166));
    InMux I__384 (
            .O(N__2191),
            .I(N__2163));
    InMux I__383 (
            .O(N__2190),
            .I(N__2152));
    InMux I__382 (
            .O(N__2189),
            .I(N__2152));
    InMux I__381 (
            .O(N__2188),
            .I(N__2152));
    InMux I__380 (
            .O(N__2187),
            .I(N__2152));
    InMux I__379 (
            .O(N__2186),
            .I(N__2152));
    CascadeMux I__378 (
            .O(N__2185),
            .I(N__2147));
    LocalMux I__377 (
            .O(N__2180),
            .I(N__2139));
    LocalMux I__376 (
            .O(N__2175),
            .I(N__2139));
    LocalMux I__375 (
            .O(N__2166),
            .I(N__2139));
    LocalMux I__374 (
            .O(N__2163),
            .I(N__2134));
    LocalMux I__373 (
            .O(N__2152),
            .I(N__2134));
    CascadeMux I__372 (
            .O(N__2151),
            .I(N__2130));
    InMux I__371 (
            .O(N__2150),
            .I(N__2125));
    InMux I__370 (
            .O(N__2147),
            .I(N__2125));
    CascadeMux I__369 (
            .O(N__2146),
            .I(N__2122));
    Span4Mux_v I__368 (
            .O(N__2139),
            .I(N__2117));
    Span4Mux_v I__367 (
            .O(N__2134),
            .I(N__2114));
    InMux I__366 (
            .O(N__2133),
            .I(N__2109));
    InMux I__365 (
            .O(N__2130),
            .I(N__2109));
    LocalMux I__364 (
            .O(N__2125),
            .I(N__2106));
    InMux I__363 (
            .O(N__2122),
            .I(N__2103));
    InMux I__362 (
            .O(N__2121),
            .I(N__2098));
    InMux I__361 (
            .O(N__2120),
            .I(N__2098));
    Odrv4 I__360 (
            .O(N__2117),
            .I(S2_S3_c_0));
    Odrv4 I__359 (
            .O(N__2114),
            .I(S2_S3_c_0));
    LocalMux I__358 (
            .O(N__2109),
            .I(S2_S3_c_0));
    Odrv4 I__357 (
            .O(N__2106),
            .I(S2_S3_c_0));
    LocalMux I__356 (
            .O(N__2103),
            .I(S2_S3_c_0));
    LocalMux I__355 (
            .O(N__2098),
            .I(S2_S3_c_0));
    CascadeMux I__354 (
            .O(N__2085),
            .I(N__2075));
    InMux I__353 (
            .O(N__2084),
            .I(N__2065));
    InMux I__352 (
            .O(N__2083),
            .I(N__2060));
    InMux I__351 (
            .O(N__2082),
            .I(N__2060));
    InMux I__350 (
            .O(N__2081),
            .I(N__2055));
    InMux I__349 (
            .O(N__2080),
            .I(N__2055));
    InMux I__348 (
            .O(N__2079),
            .I(N__2044));
    InMux I__347 (
            .O(N__2078),
            .I(N__2044));
    InMux I__346 (
            .O(N__2075),
            .I(N__2044));
    InMux I__345 (
            .O(N__2074),
            .I(N__2044));
    InMux I__344 (
            .O(N__2073),
            .I(N__2044));
    InMux I__343 (
            .O(N__2072),
            .I(N__2033));
    InMux I__342 (
            .O(N__2071),
            .I(N__2033));
    InMux I__341 (
            .O(N__2070),
            .I(N__2033));
    InMux I__340 (
            .O(N__2069),
            .I(N__2033));
    InMux I__339 (
            .O(N__2068),
            .I(N__2033));
    LocalMux I__338 (
            .O(N__2065),
            .I(N__2024));
    LocalMux I__337 (
            .O(N__2060),
            .I(N__2024));
    LocalMux I__336 (
            .O(N__2055),
            .I(N__2024));
    LocalMux I__335 (
            .O(N__2044),
            .I(N__2015));
    LocalMux I__334 (
            .O(N__2033),
            .I(N__2015));
    InMux I__333 (
            .O(N__2032),
            .I(N__2010));
    InMux I__332 (
            .O(N__2031),
            .I(N__2010));
    Span4Mux_v I__331 (
            .O(N__2024),
            .I(N__2003));
    InMux I__330 (
            .O(N__2023),
            .I(N__1994));
    InMux I__329 (
            .O(N__2022),
            .I(N__1994));
    InMux I__328 (
            .O(N__2021),
            .I(N__1994));
    InMux I__327 (
            .O(N__2020),
            .I(N__1994));
    Span4Mux_v I__326 (
            .O(N__2015),
            .I(N__1989));
    LocalMux I__325 (
            .O(N__2010),
            .I(N__1989));
    InMux I__324 (
            .O(N__2009),
            .I(N__1980));
    InMux I__323 (
            .O(N__2008),
            .I(N__1980));
    InMux I__322 (
            .O(N__2007),
            .I(N__1980));
    InMux I__321 (
            .O(N__2006),
            .I(N__1980));
    Odrv4 I__320 (
            .O(N__2003),
            .I(S2_S3_c_1));
    LocalMux I__319 (
            .O(N__1994),
            .I(S2_S3_c_1));
    Odrv4 I__318 (
            .O(N__1989),
            .I(S2_S3_c_1));
    LocalMux I__317 (
            .O(N__1980),
            .I(S2_S3_c_1));
    CascadeMux I__316 (
            .O(N__1971),
            .I(SYNTHESIZED_WIRE_0_6_cascade_));
    InMux I__315 (
            .O(N__1968),
            .I(N__1958));
    InMux I__314 (
            .O(N__1967),
            .I(N__1955));
    InMux I__313 (
            .O(N__1966),
            .I(N__1950));
    InMux I__312 (
            .O(N__1965),
            .I(N__1950));
    InMux I__311 (
            .O(N__1964),
            .I(N__1947));
    InMux I__310 (
            .O(N__1963),
            .I(N__1942));
    InMux I__309 (
            .O(N__1962),
            .I(N__1942));
    InMux I__308 (
            .O(N__1961),
            .I(N__1939));
    LocalMux I__307 (
            .O(N__1958),
            .I(N__1936));
    LocalMux I__306 (
            .O(N__1955),
            .I(N__1929));
    LocalMux I__305 (
            .O(N__1950),
            .I(N__1929));
    LocalMux I__304 (
            .O(N__1947),
            .I(N__1929));
    LocalMux I__303 (
            .O(N__1942),
            .I(N__1924));
    LocalMux I__302 (
            .O(N__1939),
            .I(N__1924));
    Span4Mux_v I__301 (
            .O(N__1936),
            .I(N__1919));
    Span4Mux_v I__300 (
            .O(N__1929),
            .I(N__1919));
    Span4Mux_v I__299 (
            .O(N__1924),
            .I(N__1916));
    Span4Mux_v I__298 (
            .O(N__1919),
            .I(N__1913));
    Span4Mux_v I__297 (
            .O(N__1916),
            .I(N__1910));
    Odrv4 I__296 (
            .O(N__1913),
            .I(S1_c));
    Odrv4 I__295 (
            .O(N__1910),
            .I(S1_c));
    InMux I__294 (
            .O(N__1905),
            .I(N__1902));
    LocalMux I__293 (
            .O(N__1902),
            .I(\b2v_inst4.result_reg2_bmZ0Z_6 ));
    InMux I__292 (
            .O(N__1899),
            .I(N__1896));
    LocalMux I__291 (
            .O(N__1896),
            .I(\b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4 ));
    InMux I__290 (
            .O(N__1893),
            .I(\b2v_inst.un8_result_arith_cry_0 ));
    InMux I__289 (
            .O(N__1890),
            .I(N__1887));
    LocalMux I__288 (
            .O(N__1887),
            .I(\b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4 ));
    InMux I__287 (
            .O(N__1884),
            .I(\b2v_inst.un8_result_arith_cry_1 ));
    InMux I__286 (
            .O(N__1881),
            .I(N__1878));
    LocalMux I__285 (
            .O(N__1878),
            .I(\b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4 ));
    InMux I__284 (
            .O(N__1875),
            .I(\b2v_inst.un8_result_arith_cry_2 ));
    InMux I__283 (
            .O(N__1872),
            .I(N__1869));
    LocalMux I__282 (
            .O(N__1869),
            .I(un8_result_arith_cry_3_c_RNIO6R4));
    InMux I__281 (
            .O(N__1866),
            .I(\b2v_inst.un8_result_arith_cry_3 ));
    InMux I__280 (
            .O(N__1863),
            .I(N__1860));
    LocalMux I__279 (
            .O(N__1860),
            .I(\b2v_inst3.result_reg1_amZ0Z_3 ));
    InMux I__278 (
            .O(N__1857),
            .I(N__1854));
    LocalMux I__277 (
            .O(N__1854),
            .I(\b2v_inst.A_equal_B_NEZ0Z_1 ));
    CascadeMux I__276 (
            .O(N__1851),
            .I(\b2v_inst3.result_reg1_bmZ0Z_2_cascade_ ));
    InMux I__275 (
            .O(N__1848),
            .I(N__1845));
    LocalMux I__274 (
            .O(N__1845),
            .I(\b2v_inst3.result_reg1_amZ0Z_2 ));
    CascadeMux I__273 (
            .O(N__1842),
            .I(SYNTHESIZED_WIRE_3_2_cascade_));
    IoInMux I__272 (
            .O(N__1839),
            .I(N__1836));
    LocalMux I__271 (
            .O(N__1836),
            .I(N__1833));
    Span4Mux_s0_h I__270 (
            .O(N__1833),
            .I(N__1830));
    Span4Mux_v I__269 (
            .O(N__1830),
            .I(N__1827));
    Odrv4 I__268 (
            .O(N__1827),
            .I(SYNTHESIZED_WIRE_4_2));
    InMux I__267 (
            .O(N__1824),
            .I(N__1821));
    LocalMux I__266 (
            .O(N__1821),
            .I(\b2v_inst.A_equal_B_NEZ0Z_3 ));
    InMux I__265 (
            .O(N__1818),
            .I(N__1815));
    LocalMux I__264 (
            .O(N__1815),
            .I(\b2v_inst.result_arith_1_2 ));
    InMux I__263 (
            .O(N__1812),
            .I(N__1809));
    LocalMux I__262 (
            .O(N__1809),
            .I(N_23));
    InMux I__261 (
            .O(N__1806),
            .I(N__1794));
    InMux I__260 (
            .O(N__1805),
            .I(N__1794));
    InMux I__259 (
            .O(N__1804),
            .I(N__1789));
    InMux I__258 (
            .O(N__1803),
            .I(N__1789));
    InMux I__257 (
            .O(N__1802),
            .I(N__1784));
    InMux I__256 (
            .O(N__1801),
            .I(N__1784));
    InMux I__255 (
            .O(N__1800),
            .I(N__1781));
    InMux I__254 (
            .O(N__1799),
            .I(N__1778));
    LocalMux I__253 (
            .O(N__1794),
            .I(N__1773));
    LocalMux I__252 (
            .O(N__1789),
            .I(N__1773));
    LocalMux I__251 (
            .O(N__1784),
            .I(N__1770));
    LocalMux I__250 (
            .O(N__1781),
            .I(N__1761));
    LocalMux I__249 (
            .O(N__1778),
            .I(N__1761));
    Sp12to4 I__248 (
            .O(N__1773),
            .I(N__1761));
    Sp12to4 I__247 (
            .O(N__1770),
            .I(N__1761));
    Span12Mux_v I__246 (
            .O(N__1761),
            .I(N__1758));
    Odrv12 I__245 (
            .O(N__1758),
            .I(s2_c));
    IoInMux I__244 (
            .O(N__1755),
            .I(N__1752));
    LocalMux I__243 (
            .O(N__1752),
            .I(N__1749));
    Odrv12 I__242 (
            .O(N__1749),
            .I(SYNTHESIZED_WIRE_4_6));
    InMux I__241 (
            .O(N__1746),
            .I(N__1743));
    LocalMux I__240 (
            .O(N__1743),
            .I(\b2v_inst.A_c_i_6 ));
    InMux I__239 (
            .O(N__1740),
            .I(N__1737));
    LocalMux I__238 (
            .O(N__1737),
            .I(\b2v_inst.A_c_i_7 ));
    InMux I__237 (
            .O(N__1734),
            .I(bfn_1_14_0_));
    IoInMux I__236 (
            .O(N__1731),
            .I(N__1727));
    CascadeMux I__235 (
            .O(N__1730),
            .I(N__1724));
    LocalMux I__234 (
            .O(N__1727),
            .I(N__1721));
    InMux I__233 (
            .O(N__1724),
            .I(N__1718));
    Span4Mux_s2_v I__232 (
            .O(N__1721),
            .I(N__1715));
    LocalMux I__231 (
            .O(N__1718),
            .I(N__1712));
    Odrv4 I__230 (
            .O(N__1715),
            .I(B_bigger_c_THRU_CO));
    Odrv4 I__229 (
            .O(N__1712),
            .I(B_bigger_c_THRU_CO));
    CascadeMux I__228 (
            .O(N__1707),
            .I(\b2v_inst3.result_reg1_amZ0Z_1_cascade_ ));
    InMux I__227 (
            .O(N__1704),
            .I(N__1701));
    LocalMux I__226 (
            .O(N__1701),
            .I(\b2v_inst3.result_reg1_bmZ0Z_1 ));
    InMux I__225 (
            .O(N__1698),
            .I(N__1695));
    LocalMux I__224 (
            .O(N__1695),
            .I(SYNTHESIZED_WIRE_3_1));
    CascadeMux I__223 (
            .O(N__1692),
            .I(\b2v_inst3.result_reg1_bmZ0Z_3_cascade_ ));
    InMux I__222 (
            .O(N__1689),
            .I(N__1686));
    LocalMux I__221 (
            .O(N__1686),
            .I(SYNTHESIZED_WIRE_3_3));
    CascadeMux I__220 (
            .O(N__1683),
            .I(N__1680));
    InMux I__219 (
            .O(N__1680),
            .I(N__1677));
    LocalMux I__218 (
            .O(N__1677),
            .I(b2v_inst_result_arith_1_7));
    InMux I__217 (
            .O(N__1674),
            .I(\b2v_inst.result_arith_1_cry_6 ));
    InMux I__216 (
            .O(N__1671),
            .I(bfn_1_12_0_));
    IoInMux I__215 (
            .O(N__1668),
            .I(N__1665));
    LocalMux I__214 (
            .O(N__1665),
            .I(N__1662));
    IoSpan4Mux I__213 (
            .O(N__1662),
            .I(N__1659));
    Sp12to4 I__212 (
            .O(N__1659),
            .I(N__1656));
    Span12Mux_s7_v I__211 (
            .O(N__1656),
            .I(N__1653));
    Odrv12 I__210 (
            .O(N__1653),
            .I(carry_out_c));
    InMux I__209 (
            .O(N__1650),
            .I(N__1647));
    LocalMux I__208 (
            .O(N__1647),
            .I(\b2v_inst.A_c_i_0 ));
    CascadeMux I__207 (
            .O(N__1644),
            .I(N__1641));
    InMux I__206 (
            .O(N__1641),
            .I(N__1638));
    LocalMux I__205 (
            .O(N__1638),
            .I(\b2v_inst.A_c_i_1 ));
    CascadeMux I__204 (
            .O(N__1635),
            .I(N__1632));
    InMux I__203 (
            .O(N__1632),
            .I(N__1629));
    LocalMux I__202 (
            .O(N__1629),
            .I(\b2v_inst.A_c_i_2 ));
    InMux I__201 (
            .O(N__1626),
            .I(N__1623));
    LocalMux I__200 (
            .O(N__1623),
            .I(\b2v_inst.A_c_i_3 ));
    InMux I__199 (
            .O(N__1620),
            .I(N__1617));
    LocalMux I__198 (
            .O(N__1617),
            .I(\b2v_inst.A_c_i_4 ));
    InMux I__197 (
            .O(N__1614),
            .I(N__1611));
    LocalMux I__196 (
            .O(N__1611),
            .I(\b2v_inst.A_c_i_5 ));
    CascadeMux I__195 (
            .O(N__1608),
            .I(\b2v_inst4.result_reg2_amZ0Z_7_cascade_ ));
    IoInMux I__194 (
            .O(N__1605),
            .I(N__1602));
    LocalMux I__193 (
            .O(N__1602),
            .I(SYNTHESIZED_WIRE_4_7));
    InMux I__192 (
            .O(N__1599),
            .I(N__1596));
    LocalMux I__191 (
            .O(N__1596),
            .I(\b2v_inst.result_arith_1_1 ));
    InMux I__190 (
            .O(N__1593),
            .I(\b2v_inst.result_arith_1_cry_0 ));
    InMux I__189 (
            .O(N__1590),
            .I(\b2v_inst.result_arith_1_cry_1 ));
    InMux I__188 (
            .O(N__1587),
            .I(N__1584));
    LocalMux I__187 (
            .O(N__1584),
            .I(\b2v_inst.result_arith_1_3 ));
    InMux I__186 (
            .O(N__1581),
            .I(\b2v_inst.result_arith_1_cry_2 ));
    CascadeMux I__185 (
            .O(N__1578),
            .I(N__1575));
    InMux I__184 (
            .O(N__1575),
            .I(N__1572));
    LocalMux I__183 (
            .O(N__1572),
            .I(b2v_inst_result_arith_1_4));
    InMux I__182 (
            .O(N__1569),
            .I(\b2v_inst.result_arith_1_cry_3 ));
    CascadeMux I__181 (
            .O(N__1566),
            .I(N__1563));
    InMux I__180 (
            .O(N__1563),
            .I(N__1560));
    LocalMux I__179 (
            .O(N__1560),
            .I(b2v_inst_result_arith_1_5));
    InMux I__178 (
            .O(N__1557),
            .I(\b2v_inst.result_arith_1_cry_4 ));
    InMux I__177 (
            .O(N__1554),
            .I(\b2v_inst.result_arith_1_cry_5 ));
    CascadeMux I__176 (
            .O(N__1551),
            .I(\b2v_inst4.result_reg2_bmZ0Z_4_cascade_ ));
    IoInMux I__175 (
            .O(N__1548),
            .I(N__1545));
    LocalMux I__174 (
            .O(N__1545),
            .I(N__1542));
    IoSpan4Mux I__173 (
            .O(N__1542),
            .I(N__1539));
    Odrv4 I__172 (
            .O(N__1539),
            .I(SYNTHESIZED_WIRE_4_4));
    CascadeMux I__171 (
            .O(N__1536),
            .I(SYNTHESIZED_WIRE_0_5_cascade_));
    CascadeMux I__170 (
            .O(N__1533),
            .I(\b2v_inst4.result_reg2_bmZ0Z_5_cascade_ ));
    IoInMux I__169 (
            .O(N__1530),
            .I(N__1527));
    LocalMux I__168 (
            .O(N__1527),
            .I(SYNTHESIZED_WIRE_4_5));
    CascadeMux I__167 (
            .O(N__1524),
            .I(N__1521));
    InMux I__166 (
            .O(N__1521),
            .I(N__1518));
    LocalMux I__165 (
            .O(N__1518),
            .I(N__1515));
    Odrv12 I__164 (
            .O(N__1515),
            .I(N_22));
    CascadeMux I__163 (
            .O(N__1512),
            .I(N_24_cascade_));
    IoInMux I__162 (
            .O(N__1509),
            .I(N__1506));
    LocalMux I__161 (
            .O(N__1506),
            .I(N__1503));
    Span4Mux_s0_h I__160 (
            .O(N__1503),
            .I(N__1500));
    Span4Mux_v I__159 (
            .O(N__1500),
            .I(N__1497));
    Odrv4 I__158 (
            .O(N__1497),
            .I(SYNTHESIZED_WIRE_4_3));
    InMux I__157 (
            .O(N__1494),
            .I(N__1491));
    LocalMux I__156 (
            .O(N__1491),
            .I(\b2v_inst4.result_reg2_amZ0Z_4 ));
    InMux I__155 (
            .O(N__1488),
            .I(N__1485));
    LocalMux I__154 (
            .O(N__1485),
            .I(\b2v_inst4.result_reg2_amZ0Z_5 ));
    IoInMux I__153 (
            .O(N__1482),
            .I(N__1479));
    LocalMux I__152 (
            .O(N__1479),
            .I(N__1476));
    Span4Mux_s0_h I__151 (
            .O(N__1476),
            .I(N__1473));
    Odrv4 I__150 (
            .O(N__1473),
            .I(SYNTHESIZED_WIRE_4_1));
    InMux I__149 (
            .O(N__1470),
            .I(N__1467));
    LocalMux I__148 (
            .O(N__1467),
            .I(\b2v_inst3.result_reg1_bmZ0Z_0 ));
    CascadeMux I__147 (
            .O(N__1464),
            .I(\b2v_inst3.result_reg1_amZ0Z_0_cascade_ ));
    CascadeMux I__146 (
            .O(N__1461),
            .I(SYNTHESIZED_WIRE_3_0_cascade_));
    InMux I__145 (
            .O(N__1458),
            .I(N__1455));
    LocalMux I__144 (
            .O(N__1455),
            .I(N_21));
    IoInMux I__143 (
            .O(N__1452),
            .I(N__1449));
    LocalMux I__142 (
            .O(N__1449),
            .I(N__1446));
    IoSpan4Mux I__141 (
            .O(N__1446),
            .I(N__1443));
    Odrv4 I__140 (
            .O(N__1443),
            .I(SYNTHESIZED_WIRE_4_0));
    CascadeMux I__139 (
            .O(N__1440),
            .I(\b2v_inst.A_equal_B_NEZ0Z_2_cascade_ ));
    InMux I__138 (
            .O(N__1437),
            .I(N__1434));
    LocalMux I__137 (
            .O(N__1434),
            .I(\b2v_inst.A_equal_B_NEZ0Z_0 ));
    IoInMux I__136 (
            .O(N__1431),
            .I(N__1428));
    LocalMux I__135 (
            .O(N__1428),
            .I(N__1425));
    IoSpan4Mux I__134 (
            .O(N__1425),
            .I(N__1422));
    IoSpan4Mux I__133 (
            .O(N__1422),
            .I(N__1419));
    Odrv4 I__132 (
            .O(N__1419),
            .I(A_equal_B_c));
    CascadeMux I__131 (
            .O(N__1416),
            .I(SYNTHESIZED_WIRE_0_4_cascade_));
    ClkMux I__130 (
            .O(N__1413),
            .I(N__1398));
    ClkMux I__129 (
            .O(N__1412),
            .I(N__1398));
    ClkMux I__128 (
            .O(N__1411),
            .I(N__1398));
    ClkMux I__127 (
            .O(N__1410),
            .I(N__1398));
    ClkMux I__126 (
            .O(N__1409),
            .I(N__1398));
    GlobalMux I__125 (
            .O(N__1398),
            .I(N__1395));
    gio2CtrlBuf I__124 (
            .O(N__1395),
            .I(CLK_c_g));
    IoInMux I__123 (
            .O(N__1392),
            .I(N__1389));
    LocalMux I__122 (
            .O(N__1389),
            .I(CONSTANT_ONE_NET));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\b2v_inst.result_arith_1_8 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(B_bigger_c),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(A_bigger_c),
            .carryinitout(bfn_2_13_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_3_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_3_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_3_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_bm_0_LC_1_8_1 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_bm_0_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_bm_0_LC_1_8_1 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \b2v_inst3.result_reg1_bm_0_LC_1_8_1  (
            .in0(N__2322),
            .in1(N__2007),
            .in2(N__2146),
            .in3(N__2667),
            .lcout(\b2v_inst3.result_reg1_bmZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_0_0_LC_1_8_2 .C_ON=1'b0;
    defparam \b2v_inst.result_arith_0_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_0_0_LC_1_8_2 .LUT_INIT=16'b0001111010110100;
    LogicCell40 \b2v_inst.result_arith_0_0_LC_1_8_2  (
            .in0(N__2120),
            .in1(N__2785),
            .in2(N__2844),
            .in3(N__2786),
            .lcout(N_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_equal_B_NE_0_LC_1_8_3 .C_ON=1'b0;
    defparam \b2v_inst.A_equal_B_NE_0_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_equal_B_NE_0_LC_1_8_3 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \b2v_inst.A_equal_B_NE_0_LC_1_8_3  (
            .in0(N__2577),
            .in1(N__2666),
            .in2(N__2843),
            .in3(N__2784),
            .lcout(\b2v_inst.A_equal_B_NEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_1_LC_1_8_4 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_1_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_1_LC_1_8_4 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \b2v_inst4.result_reg2_1_LC_1_8_4  (
            .in0(N__2009),
            .in1(N__1802),
            .in2(N__1524),
            .in3(N__1698),
            .lcout(SYNTHESIZED_WIRE_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_am_0_LC_1_8_5 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_am_0_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_am_0_LC_1_8_5 .LUT_INIT=16'b0101011001100100;
    LogicCell40 \b2v_inst3.result_reg1_am_0_LC_1_8_5  (
            .in0(N__2838),
            .in1(N__2006),
            .in2(N__2790),
            .in3(N__2121),
            .lcout(),
            .ltout(\b2v_inst3.result_reg1_amZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_ns_0_LC_1_8_6 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_ns_0_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_ns_0_LC_1_8_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \b2v_inst3.result_reg1_ns_0_LC_1_8_6  (
            .in0(N__1470),
            .in1(_gnd_net_),
            .in2(N__1464),
            .in3(N__1961),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_0_LC_1_8_7 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_0_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_0_LC_1_8_7 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \b2v_inst4.result_reg2_0_LC_1_8_7  (
            .in0(N__1801),
            .in1(N__2008),
            .in2(N__1461),
            .in3(N__1458),
            .lcout(SYNTHESIZED_WIRE_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_equal_B_NE_2_LC_1_9_0 .C_ON=1'b0;
    defparam \b2v_inst.A_equal_B_NE_2_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_equal_B_NE_2_LC_1_9_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \b2v_inst.A_equal_B_NE_2_LC_1_9_0  (
            .in0(N__3263),
            .in1(N__3217),
            .in2(N__3324),
            .in3(N__3379),
            .lcout(),
            .ltout(\b2v_inst.A_equal_B_NEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_equal_B_NE_LC_1_9_1 .C_ON=1'b0;
    defparam \b2v_inst.A_equal_B_NE_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_equal_B_NE_LC_1_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.A_equal_B_NE_LC_1_9_1  (
            .in0(N__1857),
            .in1(N__1824),
            .in2(N__1440),
            .in3(N__1437),
            .lcout(A_equal_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.result_logic_4_LC_1_9_2 .C_ON=1'b0;
    defparam \b2v_inst1.result_logic_4_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.result_logic_4_LC_1_9_2 .LUT_INIT=16'b0101011001100100;
    LogicCell40 \b2v_inst1.result_logic_4_LC_1_9_2  (
            .in0(N__3322),
            .in1(N__2020),
            .in2(N__2151),
            .in3(N__3380),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_bm_4_LC_1_9_3 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_bm_4_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_bm_4_LC_1_9_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst4.result_reg2_bm_4_LC_1_9_3  (
            .in0(N__2022),
            .in1(N__1962),
            .in2(N__1416),
            .in3(N__2324),
            .lcout(),
            .ltout(\b2v_inst4.result_reg2_bmZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_ns_4_LC_1_9_4 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_ns_4_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_ns_4_LC_1_9_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \b2v_inst4.result_reg2_ns_4_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__1803),
            .in2(N__1551),
            .in3(N__1494),
            .lcout(SYNTHESIZED_WIRE_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.result_logic_5_LC_1_9_5 .C_ON=1'b0;
    defparam \b2v_inst1.result_logic_5_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.result_logic_5_LC_1_9_5 .LUT_INIT=16'b0001010011101010;
    LogicCell40 \b2v_inst1.result_logic_5_LC_1_9_5  (
            .in0(N__2021),
            .in1(N__2133),
            .in2(N__3225),
            .in3(N__3264),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_bm_5_LC_1_9_6 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_bm_5_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_bm_5_LC_1_9_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst4.result_reg2_bm_5_LC_1_9_6  (
            .in0(N__1963),
            .in1(N__3381),
            .in2(N__1536),
            .in3(N__2023),
            .lcout(),
            .ltout(\b2v_inst4.result_reg2_bmZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_ns_5_LC_1_9_7 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_ns_5_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_ns_5_LC_1_9_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst4.result_reg2_ns_5_LC_1_9_7  (
            .in0(N__1804),
            .in1(_gnd_net_),
            .in2(N__1533),
            .in3(N__1488),
            .lcout(SYNTHESIZED_WIRE_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNI1KOT_LC_1_10_0 .C_ON=1'b0;
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNI1KOT_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNI1KOT_LC_1_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.un8_result_arith_cry_0_c_RNI1KOT_LC_1_10_0  (
            .in0(N__1599),
            .in1(N__1899),
            .in2(_gnd_net_),
            .in3(N__2186),
            .lcout(N_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIB2TT_LC_1_10_1 .C_ON=1'b0;
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIB2TT_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIB2TT_LC_1_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst.un8_result_arith_cry_2_c_RNIB2TT_LC_1_10_1  (
            .in0(N__2187),
            .in1(N__1881),
            .in2(_gnd_net_),
            .in3(N__1587),
            .lcout(),
            .ltout(N_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_3_LC_1_10_2 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_3_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_3_LC_1_10_2 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \b2v_inst4.result_reg2_3_LC_1_10_2  (
            .in0(N__1805),
            .in1(N__1689),
            .in2(N__1512),
            .in3(N__2080),
            .lcout(SYNTHESIZED_WIRE_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_am_4_LC_1_10_4 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_am_4_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_am_4_LC_1_10_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \b2v_inst4.result_reg2_am_4_LC_1_10_4  (
            .in0(N__1872),
            .in1(N__2081),
            .in2(N__1578),
            .in3(N__2188),
            .lcout(\b2v_inst4.result_reg2_amZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_am_5_LC_1_10_5 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_am_5_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_am_5_LC_1_10_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \b2v_inst4.result_reg2_am_5_LC_1_10_5  (
            .in0(N__2189),
            .in1(N__2871),
            .in2(N__1566),
            .in3(N__2082),
            .lcout(\b2v_inst4.result_reg2_amZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_am_7_LC_1_10_6 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_am_7_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_am_7_LC_1_10_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst4.result_reg2_am_7_LC_1_10_6  (
            .in0(N__2083),
            .in1(N__2850),
            .in2(N__1683),
            .in3(N__2190),
            .lcout(),
            .ltout(\b2v_inst4.result_reg2_amZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_ns_7_LC_1_10_7 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_ns_7_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_ns_7_LC_1_10_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \b2v_inst4.result_reg2_ns_7_LC_1_10_7  (
            .in0(N__2220),
            .in1(_gnd_net_),
            .in2(N__1608),
            .in3(N__1806),
            .lcout(SYNTHESIZED_WIRE_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_0_c_LC_1_11_0 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_0_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_0_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.result_arith_1_cry_0_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__2805),
            .in2(N__2782),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\b2v_inst.result_arith_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_0_c_RNIOBEO_LC_1_11_1 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_0_c_RNIOBEO_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_0_c_RNIOBEO_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_0_c_RNIOBEO_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__2549),
            .in2(N__2664),
            .in3(N__1593),
            .lcout(\b2v_inst.result_arith_1_1 ),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_0 ),
            .carryout(\b2v_inst.result_arith_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_1_c_RNIRFFO_LC_1_11_2 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_1_c_RNIRFFO_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_1_c_RNIRFFO_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_1_c_RNIRFFO_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__2515),
            .in2(N__2436),
            .in3(N__1590),
            .lcout(\b2v_inst.result_arith_1_2 ),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_1 ),
            .carryout(\b2v_inst.result_arith_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_2_c_RNIUJGO_LC_1_11_3 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_2_c_RNIUJGO_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_2_c_RNIUJGO_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_2_c_RNIUJGO_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__2379),
            .in2(N__2331),
            .in3(N__1581),
            .lcout(\b2v_inst.result_arith_1_3 ),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_2 ),
            .carryout(\b2v_inst.result_arith_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_3_c_RNI1OHO_LC_1_11_4 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_3_c_RNI1OHO_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_3_c_RNI1OHO_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_3_c_RNI1OHO_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__3306),
            .in2(N__3378),
            .in3(N__1569),
            .lcout(b2v_inst_result_arith_1_4),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_3 ),
            .carryout(\b2v_inst.result_arith_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_4_c_RNI4SIO_LC_1_11_5 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_4_c_RNI4SIO_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_4_c_RNI4SIO_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_4_c_RNI4SIO_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__3252),
            .in2(N__3222),
            .in3(N__1557),
            .lcout(b2v_inst_result_arith_1_5),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_4 ),
            .carryout(\b2v_inst.result_arith_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_5_c_RNI70KO_LC_1_11_6 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_5_c_RNI70KO_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_5_c_RNI70KO_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_5_c_RNI70KO_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__3124),
            .in2(N__3083),
            .in3(N__1554),
            .lcout(b2v_inst_result_arith_1_6),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_5 ),
            .carryout(\b2v_inst.result_arith_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_6_c_RNIA4LO_LC_1_11_7 .C_ON=1'b1;
    defparam \b2v_inst.result_arith_1_cry_6_c_RNIA4LO_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_6_c_RNIA4LO_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.result_arith_1_cry_6_c_RNIA4LO_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__2990),
            .in2(N__2947),
            .in3(N__1674),
            .lcout(b2v_inst_result_arith_1_7),
            .ltout(),
            .carryin(\b2v_inst.result_arith_1_cry_6 ),
            .carryout(\b2v_inst.result_arith_1_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.result_arith_1_cry_7_c_RNIQ27A_LC_1_12_0 .C_ON=1'b0;
    defparam \b2v_inst.result_arith_1_cry_7_c_RNIQ27A_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.result_arith_1_cry_7_c_RNIQ27A_LC_1_12_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \b2v_inst.result_arith_1_cry_7_c_RNIQ27A_LC_1_12_0  (
            .in0(N__2191),
            .in1(N__2084),
            .in2(N__1730),
            .in3(N__1671),
            .lcout(carry_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_0_c_inv_LC_1_13_0 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_0_c_inv_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_0_c_inv_LC_1_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.B_bigger_cry_0_c_inv_LC_1_13_0  (
            .in0(N__2751),
            .in1(N__1650),
            .in2(N__2842),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.A_c_i_0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\b2v_inst.B_bigger_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_1_c_inv_LC_1_13_1 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_1_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_1_c_inv_LC_1_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.B_bigger_cry_1_c_inv_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__2576),
            .in2(N__1644),
            .in3(N__2643),
            .lcout(\b2v_inst.A_c_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_0 ),
            .carryout(\b2v_inst.B_bigger_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_2_c_inv_LC_1_13_2 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_2_c_inv_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_2_c_inv_LC_1_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.B_bigger_cry_2_c_inv_LC_1_13_2  (
            .in0(N__2501),
            .in1(N__2421),
            .in2(N__1635),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.A_c_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_1 ),
            .carryout(\b2v_inst.B_bigger_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_3_c_inv_LC_1_13_3 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_3_c_inv_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_3_c_inv_LC_1_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.B_bigger_cry_3_c_inv_LC_1_13_3  (
            .in0(N__2287),
            .in1(N__1626),
            .in2(N__2378),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.A_c_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_2 ),
            .carryout(\b2v_inst.B_bigger_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_4_c_inv_LC_1_13_4 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_4_c_inv_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_4_c_inv_LC_1_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.B_bigger_cry_4_c_inv_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__1620),
            .in2(N__3323),
            .in3(N__3340),
            .lcout(\b2v_inst.A_c_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_3 ),
            .carryout(\b2v_inst.B_bigger_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_5_c_inv_LC_1_13_5 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_5_c_inv_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_5_c_inv_LC_1_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.B_bigger_cry_5_c_inv_LC_1_13_5  (
            .in0(N__3199),
            .in1(N__1614),
            .in2(N__3257),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.A_c_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_4 ),
            .carryout(\b2v_inst.B_bigger_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_6_c_inv_LC_1_13_6 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_6_c_inv_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_6_c_inv_LC_1_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.B_bigger_cry_6_c_inv_LC_1_13_6  (
            .in0(N__3043),
            .in1(N__1746),
            .in2(N__3111),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.A_c_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_5 ),
            .carryout(\b2v_inst.B_bigger_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.B_bigger_cry_7_c_inv_LC_1_13_7 .C_ON=1'b1;
    defparam \b2v_inst.B_bigger_cry_7_c_inv_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.B_bigger_cry_7_c_inv_LC_1_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.B_bigger_cry_7_c_inv_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__1740),
            .in2(N__3000),
            .in3(N__2910),
            .lcout(\b2v_inst.A_c_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.B_bigger_cry_6 ),
            .carryout(B_bigger_c),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_bigger_c_THRU_LUT4_0_LC_1_14_0.C_ON=1'b0;
    defparam B_bigger_c_THRU_LUT4_0_LC_1_14_0.SEQ_MODE=4'b0000;
    defparam B_bigger_c_THRU_LUT4_0_LC_1_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 B_bigger_c_THRU_LUT4_0_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1734),
            .lcout(B_bigger_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_bm_1_LC_2_8_0 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_bm_1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_bm_1_LC_2_8_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \b2v_inst3.result_reg1_bm_1_LC_2_8_0  (
            .in0(N__2771),
            .in1(N__2032),
            .in2(N__2516),
            .in3(N__2150),
            .lcout(\b2v_inst3.result_reg1_bmZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_am_1_LC_2_8_1 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_am_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_am_1_LC_2_8_1 .LUT_INIT=16'b0001010011101010;
    LogicCell40 \b2v_inst3.result_reg1_am_1_LC_2_8_1  (
            .in0(N__2031),
            .in1(N__2657),
            .in2(N__2185),
            .in3(N__2575),
            .lcout(),
            .ltout(\b2v_inst3.result_reg1_amZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_ns_1_LC_2_8_2 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_ns_1_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_ns_1_LC_2_8_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst3.result_reg1_ns_1_LC_2_8_2  (
            .in0(N__1964),
            .in1(_gnd_net_),
            .in2(N__1707),
            .in3(N__1704),
            .lcout(SYNTHESIZED_WIRE_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_bm_3_LC_2_9_0 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_bm_3_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_bm_3_LC_2_9_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \b2v_inst3.result_reg1_bm_3_LC_2_9_0  (
            .in0(N__2195),
            .in1(N__2071),
            .in2(N__2783),
            .in3(N__2494),
            .lcout(),
            .ltout(\b2v_inst3.result_reg1_bmZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_ns_3_LC_2_9_1 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_ns_3_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_ns_3_LC_2_9_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst3.result_reg1_ns_3_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__1863),
            .in2(N__1692),
            .in3(N__1966),
            .lcout(SYNTHESIZED_WIRE_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_am_2_LC_2_9_2 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_am_2_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_am_2_LC_2_9_2 .LUT_INIT=16'b0001111000101100;
    LogicCell40 \b2v_inst3.result_reg1_am_2_LC_2_9_2  (
            .in0(N__2192),
            .in1(N__2068),
            .in2(N__2448),
            .in3(N__2493),
            .lcout(\b2v_inst3.result_reg1_amZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_am_3_LC_2_9_3 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_am_3_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_am_3_LC_2_9_3 .LUT_INIT=16'b0001111001001010;
    LogicCell40 \b2v_inst3.result_reg1_am_3_LC_2_9_3  (
            .in0(N__2069),
            .in1(N__2193),
            .in2(N__2377),
            .in3(N__2329),
            .lcout(\b2v_inst3.result_reg1_amZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_equal_B_NE_1_LC_2_9_4 .C_ON=1'b0;
    defparam \b2v_inst.A_equal_B_NE_1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_equal_B_NE_1_LC_2_9_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \b2v_inst.A_equal_B_NE_1_LC_2_9_4  (
            .in0(N__2328),
            .in1(N__2367),
            .in2(N__2447),
            .in3(N__2492),
            .lcout(\b2v_inst.A_equal_B_NEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_bm_2_LC_2_9_5 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_bm_2_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_bm_2_LC_2_9_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \b2v_inst3.result_reg1_bm_2_LC_2_9_5  (
            .in0(N__2070),
            .in1(N__2330),
            .in2(N__2665),
            .in3(N__2194),
            .lcout(),
            .ltout(\b2v_inst3.result_reg1_bmZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.result_reg1_ns_2_LC_2_9_6 .C_ON=1'b0;
    defparam \b2v_inst3.result_reg1_ns_2_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.result_reg1_ns_2_LC_2_9_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst3.result_reg1_ns_2_LC_2_9_6  (
            .in0(N__1965),
            .in1(_gnd_net_),
            .in2(N__1851),
            .in3(N__1848),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_3_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_2_LC_2_9_7 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_2_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_2_LC_2_9_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \b2v_inst4.result_reg2_2_LC_2_9_7  (
            .in0(N__2072),
            .in1(N__1812),
            .in2(N__1842),
            .in3(N__1799),
            .lcout(SYNTHESIZED_WIRE_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_equal_B_NE_3_LC_2_10_0 .C_ON=1'b0;
    defparam \b2v_inst.A_equal_B_NE_3_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_equal_B_NE_3_LC_2_10_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \b2v_inst.A_equal_B_NE_3_LC_2_10_0  (
            .in0(N__3014),
            .in1(N__3125),
            .in2(N__3090),
            .in3(N__2948),
            .lcout(\b2v_inst.A_equal_B_NEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNI6RQT_LC_2_10_1 .C_ON=1'b0;
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNI6RQT_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNI6RQT_LC_2_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst.un8_result_arith_cry_1_c_RNI6RQT_LC_2_10_1  (
            .in0(N__2196),
            .in1(N__1890),
            .in2(_gnd_net_),
            .in3(N__1818),
            .lcout(N_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_ns_6_LC_2_10_2 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_ns_6_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_ns_6_LC_2_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst4.result_reg2_ns_6_LC_2_10_2  (
            .in0(N__2208),
            .in1(N__1800),
            .in2(_gnd_net_),
            .in3(N__1905),
            .lcout(SYNTHESIZED_WIRE_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.result_logic_7_LC_2_10_3 .C_ON=1'b0;
    defparam \b2v_inst1.result_logic_7_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.result_logic_7_LC_2_10_3 .LUT_INIT=16'b0001010011101010;
    LogicCell40 \b2v_inst1.result_logic_7_LC_2_10_3  (
            .in0(N__2074),
            .in1(N__2201),
            .in2(N__2952),
            .in3(N__3015),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_bm_7_LC_2_10_4 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_bm_7_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_bm_7_LC_2_10_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst4.result_reg2_bm_7_LC_2_10_4  (
            .in0(N__3089),
            .in1(N__2079),
            .in2(N__2223),
            .in3(N__1968),
            .lcout(\b2v_inst4.result_reg2_bmZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_am_6_LC_2_10_5 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_am_6_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_am_6_LC_2_10_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \b2v_inst4.result_reg2_am_6_LC_2_10_5  (
            .in0(N__2197),
            .in1(N__2862),
            .in2(N__2085),
            .in3(N__2214),
            .lcout(\b2v_inst4.result_reg2_amZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.result_logic_6_LC_2_10_6 .C_ON=1'b0;
    defparam \b2v_inst1.result_logic_6_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.result_logic_6_LC_2_10_6 .LUT_INIT=16'b0001001011101100;
    LogicCell40 \b2v_inst1.result_logic_6_LC_2_10_6  (
            .in0(N__3088),
            .in1(N__2073),
            .in2(N__2202),
            .in3(N__3126),
            .lcout(),
            .ltout(SYNTHESIZED_WIRE_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.result_reg2_bm_6_LC_2_10_7 .C_ON=1'b0;
    defparam \b2v_inst4.result_reg2_bm_6_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.result_reg2_bm_6_LC_2_10_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst4.result_reg2_bm_6_LC_2_10_7  (
            .in0(N__2078),
            .in1(N__3223),
            .in2(N__1971),
            .in3(N__1967),
            .lcout(\b2v_inst4.result_reg2_bmZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_0_c_LC_2_11_0 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_0_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_0_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un8_result_arith_cry_0_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__2681),
            .in2(N__2770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\b2v_inst.un8_result_arith_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNIITN4_LC_2_11_1 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNIITN4_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_0_c_RNIITN4_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_0_c_RNIITN4_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__2529),
            .in2(N__2663),
            .in3(N__1893),
            .lcout(\b2v_inst.un8_result_arith_cry_0_c_RNIITNZ0Z4 ),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_0 ),
            .carryout(\b2v_inst.un8_result_arith_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNIK0P4_LC_2_11_2 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNIK0P4_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_1_c_RNIK0P4_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_1_c_RNIK0P4_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__2391),
            .in2(N__2517),
            .in3(N__1884),
            .lcout(\b2v_inst.un8_result_arith_cry_1_c_RNIK0PZ0Z4 ),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_1 ),
            .carryout(\b2v_inst.un8_result_arith_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIM3Q4_LC_2_11_3 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIM3Q4_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_2_c_RNIM3Q4_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_2_c_RNIM3Q4_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__2235),
            .in2(N__2323),
            .in3(N__1875),
            .lcout(\b2v_inst.un8_result_arith_cry_2_c_RNIM3QZ0Z4 ),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_2 ),
            .carryout(\b2v_inst.un8_result_arith_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_3_c_RNIO6R4_LC_2_11_4 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_3_c_RNIO6R4_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_3_c_RNIO6R4_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_3_c_RNIO6R4_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__3369),
            .in2(N__3279),
            .in3(N__1866),
            .lcout(un8_result_arith_cry_3_c_RNIO6R4),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_3 ),
            .carryout(\b2v_inst.un8_result_arith_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_4_c_RNIQ9S4_LC_2_11_5 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_4_c_RNIQ9S4_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_4_c_RNIQ9S4_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_4_c_RNIQ9S4_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__3138),
            .in2(N__3221),
            .in3(N__2865),
            .lcout(un8_result_arith_cry_4_c_RNIQ9S4),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_4 ),
            .carryout(\b2v_inst.un8_result_arith_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_5_c_RNISCT4_LC_2_11_6 .C_ON=1'b1;
    defparam \b2v_inst.un8_result_arith_cry_5_c_RNISCT4_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_5_c_RNISCT4_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_result_arith_cry_5_c_RNISCT4_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__3027),
            .in2(N__3084),
            .in3(N__2856),
            .lcout(un8_result_arith_cry_5_c_RNISCT4),
            .ltout(),
            .carryin(\b2v_inst.un8_result_arith_cry_5 ),
            .carryout(\b2v_inst.un8_result_arith_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_result_arith_cry_6_c_RNIK5GH_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst.un8_result_arith_cry_6_c_RNIK5GH_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_result_arith_cry_6_c_RNIK5GH_LC_2_11_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \b2v_inst.un8_result_arith_cry_6_c_RNIK5GH_LC_2_11_7  (
            .in0(N__3012),
            .in1(N__2937),
            .in2(_gnd_net_),
            .in3(N__2853),
            .lcout(un8_result_arith_cry_6_c_RNIK5GH),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_0_c_inv_LC_2_12_0 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_0_c_inv_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_0_c_inv_LC_2_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.A_bigger_cry_0_c_inv_LC_2_12_0  (
            .in0(N__2831),
            .in1(N__2744),
            .in2(N__2682),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.B_c_i_0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\b2v_inst.A_bigger_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_1_c_inv_LC_2_12_1 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_1_c_inv_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_1_c_inv_LC_2_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.A_bigger_cry_1_c_inv_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__2528),
            .in2(N__2650),
            .in3(N__2574),
            .lcout(\b2v_inst.B_c_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_0 ),
            .carryout(\b2v_inst.A_bigger_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_2_c_inv_LC_2_12_2 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_2_c_inv_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_2_c_inv_LC_2_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.A_bigger_cry_2_c_inv_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__2390),
            .in2(N__2511),
            .in3(N__2446),
            .lcout(\b2v_inst.B_c_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_1 ),
            .carryout(\b2v_inst.A_bigger_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_3_c_inv_LC_2_12_3 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_3_c_inv_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_3_c_inv_LC_2_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.A_bigger_cry_3_c_inv_LC_2_12_3  (
            .in0(N__2360),
            .in1(N__2234),
            .in2(N__2311),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.B_c_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_2 ),
            .carryout(\b2v_inst.A_bigger_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_4_c_inv_LC_2_12_4 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_4_c_inv_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_4_c_inv_LC_2_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.A_bigger_cry_4_c_inv_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__3275),
            .in2(N__3377),
            .in3(N__3307),
            .lcout(\b2v_inst.B_c_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_3 ),
            .carryout(\b2v_inst.A_bigger_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_5_c_inv_LC_2_12_5 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_5_c_inv_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_5_c_inv_LC_2_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.A_bigger_cry_5_c_inv_LC_2_12_5  (
            .in0(N__3256),
            .in1(N__3137),
            .in2(N__3224),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.B_c_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_4 ),
            .carryout(\b2v_inst.A_bigger_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_6_c_inv_LC_2_12_6 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_6_c_inv_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_6_c_inv_LC_2_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.A_bigger_cry_6_c_inv_LC_2_12_6  (
            .in0(N__3123),
            .in1(N__3026),
            .in2(N__3082),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.B_c_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_5 ),
            .carryout(\b2v_inst.A_bigger_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.A_bigger_cry_7_c_inv_LC_2_12_7 .C_ON=1'b1;
    defparam \b2v_inst.A_bigger_cry_7_c_inv_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.A_bigger_cry_7_c_inv_LC_2_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.A_bigger_cry_7_c_inv_LC_2_12_7  (
            .in0(N__3013),
            .in1(N__2892),
            .in2(N__2946),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.B_c_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.A_bigger_cry_6 ),
            .carryout(A_bigger_c),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam A_bigger_c_THRU_LUT4_0_LC_2_13_0.C_ON=1'b0;
    defparam A_bigger_c_THRU_LUT4_0_LC_2_13_0.SEQ_MODE=4'b0000;
    defparam A_bigger_c_THRU_LUT4_0_LC_2_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 A_bigger_c_THRU_LUT4_0_LC_2_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2886),
            .lcout(A_bigger_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // ALU_STURCTURE
