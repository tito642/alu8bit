// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 22 2023 21:20:02

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "alu_behavioral" view "INTERFACE"

module alu_behavioral (
    alu_out,
    s,
    A,
    B,
    clk);

    output [7:0] alu_out;
    input [3:0] s;
    input [7:0] A;
    input [7:0] B;
    input clk;

    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2957;
    wire N__2956;
    wire N__2955;
    wire N__2948;
    wire N__2947;
    wire N__2946;
    wire N__2939;
    wire N__2938;
    wire N__2937;
    wire N__2930;
    wire N__2929;
    wire N__2928;
    wire N__2921;
    wire N__2920;
    wire N__2919;
    wire N__2912;
    wire N__2911;
    wire N__2910;
    wire N__2903;
    wire N__2902;
    wire N__2901;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2885;
    wire N__2884;
    wire N__2883;
    wire N__2876;
    wire N__2875;
    wire N__2874;
    wire N__2867;
    wire N__2866;
    wire N__2865;
    wire N__2858;
    wire N__2857;
    wire N__2856;
    wire N__2849;
    wire N__2848;
    wire N__2847;
    wire N__2840;
    wire N__2839;
    wire N__2838;
    wire N__2831;
    wire N__2830;
    wire N__2829;
    wire N__2822;
    wire N__2821;
    wire N__2820;
    wire N__2813;
    wire N__2812;
    wire N__2811;
    wire N__2804;
    wire N__2803;
    wire N__2802;
    wire N__2795;
    wire N__2794;
    wire N__2793;
    wire N__2786;
    wire N__2785;
    wire N__2784;
    wire N__2777;
    wire N__2776;
    wire N__2775;
    wire N__2768;
    wire N__2767;
    wire N__2766;
    wire N__2759;
    wire N__2758;
    wire N__2757;
    wire N__2750;
    wire N__2749;
    wire N__2748;
    wire N__2741;
    wire N__2740;
    wire N__2739;
    wire N__2732;
    wire N__2731;
    wire N__2730;
    wire N__2723;
    wire N__2722;
    wire N__2721;
    wire N__2714;
    wire N__2713;
    wire N__2712;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2652;
    wire N__2647;
    wire N__2644;
    wire N__2643;
    wire N__2642;
    wire N__2637;
    wire N__2634;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2592;
    wire N__2591;
    wire N__2588;
    wire N__2581;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2569;
    wire N__2568;
    wire N__2567;
    wire N__2564;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2529;
    wire N__2528;
    wire N__2525;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2488;
    wire N__2487;
    wire N__2486;
    wire N__2485;
    wire N__2484;
    wire N__2483;
    wire N__2482;
    wire N__2481;
    wire N__2480;
    wire N__2479;
    wire N__2478;
    wire N__2469;
    wire N__2466;
    wire N__2459;
    wire N__2452;
    wire N__2451;
    wire N__2446;
    wire N__2441;
    wire N__2440;
    wire N__2439;
    wire N__2438;
    wire N__2437;
    wire N__2434;
    wire N__2433;
    wire N__2432;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2418;
    wire N__2411;
    wire N__2406;
    wire N__2399;
    wire N__2392;
    wire N__2391;
    wire N__2390;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2382;
    wire N__2381;
    wire N__2380;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2375;
    wire N__2374;
    wire N__2373;
    wire N__2372;
    wire N__2371;
    wire N__2368;
    wire N__2367;
    wire N__2366;
    wire N__2365;
    wire N__2364;
    wire N__2363;
    wire N__2362;
    wire N__2361;
    wire N__2352;
    wire N__2347;
    wire N__2338;
    wire N__2327;
    wire N__2318;
    wire N__2309;
    wire N__2308;
    wire N__2307;
    wire N__2304;
    wire N__2297;
    wire N__2292;
    wire N__2291;
    wire N__2290;
    wire N__2289;
    wire N__2288;
    wire N__2287;
    wire N__2286;
    wire N__2285;
    wire N__2284;
    wire N__2283;
    wire N__2280;
    wire N__2279;
    wire N__2278;
    wire N__2275;
    wire N__2268;
    wire N__2259;
    wire N__2246;
    wire N__2239;
    wire N__2230;
    wire N__2229;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2211;
    wire N__2208;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2192;
    wire N__2189;
    wire N__2184;
    wire N__2179;
    wire N__2174;
    wire N__2169;
    wire N__2168;
    wire N__2167;
    wire N__2166;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2150;
    wire N__2143;
    wire N__2140;
    wire N__2137;
    wire N__2134;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2122;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2106;
    wire N__2103;
    wire N__2098;
    wire N__2097;
    wire N__2094;
    wire N__2091;
    wire N__2086;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2071;
    wire N__2070;
    wire N__2067;
    wire N__2064;
    wire N__2063;
    wire N__2060;
    wire N__2055;
    wire N__2050;
    wire N__2047;
    wire N__2044;
    wire N__2041;
    wire N__2040;
    wire N__2039;
    wire N__2038;
    wire N__2035;
    wire N__2034;
    wire N__2033;
    wire N__2032;
    wire N__2027;
    wire N__2026;
    wire N__2025;
    wire N__2022;
    wire N__2021;
    wire N__2020;
    wire N__2019;
    wire N__2016;
    wire N__2009;
    wire N__2006;
    wire N__2001;
    wire N__1994;
    wire N__1991;
    wire N__1978;
    wire N__1975;
    wire N__1974;
    wire N__1971;
    wire N__1968;
    wire N__1965;
    wire N__1962;
    wire N__1961;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1949;
    wire N__1942;
    wire N__1939;
    wire N__1938;
    wire N__1935;
    wire N__1934;
    wire N__1933;
    wire N__1930;
    wire N__1927;
    wire N__1924;
    wire N__1919;
    wire N__1912;
    wire N__1909;
    wire N__1906;
    wire N__1903;
    wire N__1900;
    wire N__1897;
    wire N__1894;
    wire N__1891;
    wire N__1888;
    wire N__1885;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1870;
    wire N__1867;
    wire N__1864;
    wire N__1861;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1849;
    wire N__1846;
    wire N__1843;
    wire N__1840;
    wire N__1837;
    wire N__1834;
    wire N__1831;
    wire N__1828;
    wire N__1825;
    wire N__1822;
    wire N__1819;
    wire N__1816;
    wire N__1813;
    wire N__1810;
    wire N__1807;
    wire N__1804;
    wire N__1801;
    wire N__1798;
    wire N__1795;
    wire N__1792;
    wire N__1789;
    wire N__1786;
    wire N__1783;
    wire N__1782;
    wire N__1781;
    wire N__1780;
    wire N__1779;
    wire N__1778;
    wire N__1777;
    wire N__1774;
    wire N__1769;
    wire N__1760;
    wire N__1755;
    wire N__1752;
    wire N__1751;
    wire N__1750;
    wire N__1749;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1739;
    wire N__1732;
    wire N__1723;
    wire N__1720;
    wire N__1717;
    wire N__1714;
    wire N__1711;
    wire N__1708;
    wire N__1705;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1693;
    wire N__1690;
    wire N__1687;
    wire N__1684;
    wire N__1681;
    wire N__1678;
    wire N__1675;
    wire N__1672;
    wire N__1669;
    wire N__1668;
    wire N__1667;
    wire N__1666;
    wire N__1661;
    wire N__1656;
    wire N__1651;
    wire N__1648;
    wire N__1645;
    wire N__1642;
    wire N__1641;
    wire N__1640;
    wire N__1639;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1621;
    wire N__1618;
    wire N__1615;
    wire N__1612;
    wire N__1609;
    wire N__1606;
    wire N__1603;
    wire N__1600;
    wire N__1597;
    wire N__1594;
    wire N__1591;
    wire N__1588;
    wire N__1585;
    wire N__1584;
    wire N__1581;
    wire N__1578;
    wire N__1573;
    wire N__1570;
    wire N__1567;
    wire N__1564;
    wire N__1561;
    wire N__1558;
    wire N__1555;
    wire N__1552;
    wire N__1549;
    wire N__1546;
    wire N__1545;
    wire N__1540;
    wire N__1539;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1522;
    wire N__1519;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1507;
    wire N__1504;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1496;
    wire N__1495;
    wire N__1492;
    wire N__1489;
    wire N__1484;
    wire N__1477;
    wire N__1474;
    wire N__1471;
    wire N__1468;
    wire N__1465;
    wire N__1462;
    wire N__1459;
    wire N__1456;
    wire N__1453;
    wire N__1450;
    wire N__1447;
    wire N__1444;
    wire N__1441;
    wire N__1440;
    wire N__1437;
    wire N__1434;
    wire N__1433;
    wire N__1426;
    wire N__1423;
    wire N__1420;
    wire N__1417;
    wire N__1414;
    wire N__1411;
    wire N__1408;
    wire N__1405;
    wire N__1404;
    wire N__1403;
    wire N__1398;
    wire N__1395;
    wire N__1392;
    wire N__1389;
    wire N__1384;
    wire N__1381;
    wire N__1378;
    wire N__1375;
    wire N__1372;
    wire N__1369;
    wire N__1366;
    wire N__1363;
    wire N__1360;
    wire N__1357;
    wire N__1354;
    wire N__1351;
    wire N__1348;
    wire N__1345;
    wire N__1342;
    wire N__1339;
    wire N__1336;
    wire N__1333;
    wire N__1330;
    wire N__1327;
    wire N__1324;
    wire N__1321;
    wire N__1318;
    wire N__1315;
    wire N__1312;
    wire N__1309;
    wire N__1306;
    wire N__1303;
    wire N__1300;
    wire N__1297;
    wire N__1296;
    wire N__1293;
    wire N__1292;
    wire N__1291;
    wire N__1288;
    wire N__1285;
    wire N__1282;
    wire N__1279;
    wire N__1276;
    wire N__1271;
    wire N__1268;
    wire N__1267;
    wire N__1264;
    wire N__1261;
    wire N__1258;
    wire N__1255;
    wire N__1246;
    wire N__1243;
    wire N__1240;
    wire N__1237;
    wire N__1234;
    wire N__1231;
    wire N__1228;
    wire N__1225;
    wire N__1224;
    wire N__1223;
    wire N__1222;
    wire N__1221;
    wire N__1210;
    wire N__1207;
    wire N__1204;
    wire GNDG0;
    wire VCCG0;
    wire clk_c_g;
    wire alu_out_RNO_2Z0Z_1_cascade_;
    wire N_143_cascade_;
    wire alu_out_13_1;
    wire alu_out38_cascade_;
    wire un1_alu_out43_1_3_cascade_;
    wire un1_alu_out43_1_i;
    wire un1_alu_out43_1_2;
    wire alu_out40_0;
    wire N_90_cascade_;
    wire alu_out_RNO_3Z0Z_1;
    wire alu_out_13_5;
    wire N_87_cascade_;
    wire alu_out_13_4;
    wire alu_out_13_0;
    wire alu_out_13_6;
    wire s_c_i_1_cascade_;
    wire N_88;
    wire un1_A_1_cascade_;
    wire B_c_0;
    wire alu_out_RNO_2Z0Z_0_cascade_;
    wire N_142;
    wire alu_out_RNO_3Z0Z_0;
    wire B_c_1;
    wire N_85_cascade_;
    wire B_c_4;
    wire alu_out_RNO_3Z0Z_4;
    wire alu_out_RNO_2Z0Z_4_cascade_;
    wire N_146;
    wire A_c_4;
    wire alu_out_RNO_2Z0Z_5_cascade_;
    wire alu_out_RNO_3Z0Z_5;
    wire N_147;
    wire alu_out_RNO_2Z0Z_3_cascade_;
    wire alu_out_RNO_3Z0Z_3;
    wire N_145_cascade_;
    wire alu_out_13_3;
    wire A_c_2;
    wire A_c_1;
    wire alu_out_RNO_3Z0Z_2_cascade_;
    wire alu_out_RNO_2Z0Z_2;
    wire N_144_cascade_;
    wire alu_out_13_2;
    wire s_ibuf_RNI1HJVZ0Z_0;
    wire bfn_2_10_0_;
    wire un1_A_1;
    wire B_ibuf_RNIE5VR2Z0Z_0;
    wire alu_out_RNO_1Z0Z_0;
    wire un1_A_1_cry_0_c_THRU_CO;
    wire B_ibuf_RNIH05C1Z0Z_1;
    wire B_ibuf_RNI08QF1Z0Z_1;
    wire alu_out_RNO_1Z0Z_1;
    wire un1_A_1_cry_0;
    wire B_ibuf_RNI2AQF1Z0Z_2;
    wire alu_out_RNO_1Z0Z_2;
    wire un1_A_1_cry_1;
    wire B_ibuf_RNIJ25C1Z0Z_3;
    wire alu_out_RNO_1Z0Z_3;
    wire un1_A_1_cry_2;
    wire B_ibuf_RNIK35C1Z0Z_4;
    wire B_ibuf_RNI6EQF1Z0Z_4;
    wire alu_out_RNO_1Z0Z_4;
    wire un1_A_1_cry_3;
    wire B_ibuf_RNI8GQF1Z0Z_5;
    wire alu_out_RNO_1Z0Z_5;
    wire un1_A_1_cry_4;
    wire B_ibuf_RNIM55C1Z0Z_6;
    wire alu_out_RNO_1Z0Z_6;
    wire un1_A_1_cry_5;
    wire un1_A_1_cry_6;
    wire s_c_3;
    wire bfn_2_11_0_;
    wire alu_out_13_7;
    wire un1_A_1_axb_7;
    wire alu_out_RNO_3Z0Z_7;
    wire N_91;
    wire B_ibuf_RNII15C1Z0Z_2;
    wire B_c_2;
    wire N_86;
    wire B_c_5;
    wire N_89_cascade_;
    wire B_ibuf_RNIL45C1Z0Z_5;
    wire s_c_i_1;
    wire A_c_0;
    wire A_c_5;
    wire alu_out_RNO_2Z0Z_6_cascade_;
    wire alu_out_RNO_3Z0Z_6;
    wire N_148;
    wire B_c_3;
    wire A_c_3;
    wire B_ibuf_RNI4CQF1Z0Z_3;
    wire A_c_6;
    wire B_c_6;
    wire B_ibuf_RNIAIQF1Z0Z_6;
    wire A_c_7;
    wire s_c_1;
    wire s_c_0;
    wire B_c_7;
    wire s_c_2;
    wire alu_out_RNO_5Z0Z_7;
    wire alu_out_RNO_4Z0Z_7_cascade_;
    wire N_149;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2966),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__2968),
            .DIN(N__2967),
            .DOUT(N__2966),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__2968),
            .PADOUT(N__2967),
            .PADIN(N__2966),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__2957),
            .DIN(N__2956),
            .DOUT(N__2955),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__2957),
            .PADOUT(N__2956),
            .PADIN(N__2955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_7_iopad (
            .OE(N__2948),
            .DIN(N__2947),
            .DOUT(N__2946),
            .PACKAGEPIN(B[7]));
    defparam B_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_7_preio (
            .PADOEN(N__2948),
            .PADOUT(N__2947),
            .PADIN(N__2946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_6_iopad (
            .OE(N__2939),
            .DIN(N__2938),
            .DOUT(N__2937),
            .PACKAGEPIN(alu_out[6]));
    defparam alu_out_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_6_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_6_preio (
            .PADOEN(N__2939),
            .PADOUT(N__2938),
            .PADIN(N__2937),
            .CLOCKENABLE(N__1292),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1336),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1223));
    IO_PAD s_ibuf_0_iopad (
            .OE(N__2930),
            .DIN(N__2929),
            .DOUT(N__2928),
            .PACKAGEPIN(s[0]));
    defparam s_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam s_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO s_ibuf_0_preio (
            .PADOEN(N__2930),
            .PADOUT(N__2929),
            .PADIN(N__2928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(s_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__2921),
            .DIN(N__2920),
            .DOUT(N__2919),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__2921),
            .PADOUT(N__2920),
            .PADIN(N__2919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_3_iopad (
            .OE(N__2912),
            .DIN(N__2911),
            .DOUT(N__2910),
            .PACKAGEPIN(B[3]));
    defparam B_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_3_preio (
            .PADOEN(N__2912),
            .PADOUT(N__2911),
            .PADIN(N__2910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_3_iopad (
            .OE(N__2903),
            .DIN(N__2902),
            .DOUT(N__2901),
            .PACKAGEPIN(alu_out[3]));
    defparam alu_out_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_3_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_3_preio (
            .PADOEN(N__2903),
            .PADOUT(N__2902),
            .PADIN(N__2901),
            .CLOCKENABLE(N__1291),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1684),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1222));
    IO_PAD A_ibuf_3_iopad (
            .OE(N__2894),
            .DIN(N__2893),
            .DOUT(N__2892),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__2894),
            .PADOUT(N__2893),
            .PADIN(N__2892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_6_iopad (
            .OE(N__2885),
            .DIN(N__2884),
            .DOUT(N__2883),
            .PACKAGEPIN(B[6]));
    defparam B_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_6_preio (
            .PADOEN(N__2885),
            .PADOUT(N__2884),
            .PADIN(N__2883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_7_iopad (
            .OE(N__2876),
            .DIN(N__2875),
            .DOUT(N__2874),
            .PACKAGEPIN(alu_out[7]));
    defparam alu_out_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_7_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_7_preio (
            .PADOEN(N__2876),
            .PADOUT(N__2875),
            .PADIN(N__2874),
            .CLOCKENABLE(N__1291),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1720),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1222));
    IO_PAD s_ibuf_1_iopad (
            .OE(N__2867),
            .DIN(N__2866),
            .DOUT(N__2865),
            .PACKAGEPIN(s[1]));
    defparam s_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam s_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO s_ibuf_1_preio (
            .PADOEN(N__2867),
            .PADOUT(N__2866),
            .PADIN(N__2865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(s_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__2858),
            .DIN(N__2857),
            .DOUT(N__2856),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__2858),
            .PADOUT(N__2857),
            .PADIN(N__2856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_2_iopad (
            .OE(N__2849),
            .DIN(N__2848),
            .DOUT(N__2847),
            .PACKAGEPIN(B[2]));
    defparam B_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_2_preio (
            .PADOEN(N__2849),
            .PADOUT(N__2848),
            .PADIN(N__2847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_0_iopad (
            .OE(N__2840),
            .DIN(N__2839),
            .DOUT(N__2838),
            .PACKAGEPIN(alu_out[0]));
    defparam alu_out_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_0_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_0_preio (
            .PADOEN(N__2840),
            .PADOUT(N__2839),
            .PADIN(N__2838),
            .CLOCKENABLE(N__1296),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1224));
    IO_PAD A_ibuf_5_iopad (
            .OE(N__2831),
            .DIN(N__2830),
            .DOUT(N__2829),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__2831),
            .PADOUT(N__2830),
            .PADIN(N__2829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_0_iopad (
            .OE(N__2822),
            .DIN(N__2821),
            .DOUT(N__2820),
            .PACKAGEPIN(B[0]));
    defparam B_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_0_preio (
            .PADOEN(N__2822),
            .PADOUT(N__2821),
            .PADIN(N__2820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_2_iopad (
            .OE(N__2813),
            .DIN(N__2812),
            .DOUT(N__2811),
            .PACKAGEPIN(alu_out[2]));
    defparam alu_out_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_2_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_2_preio (
            .PADOEN(N__2813),
            .PADOUT(N__2812),
            .PADIN(N__2811),
            .CLOCKENABLE(N__1296),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1224));
    IO_PAD alu_out_obuf_4_iopad (
            .OE(N__2804),
            .DIN(N__2803),
            .DOUT(N__2802),
            .PACKAGEPIN(alu_out[4]));
    defparam alu_out_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_4_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_4_preio (
            .PADOEN(N__2804),
            .PADOUT(N__2803),
            .PADIN(N__2802),
            .CLOCKENABLE(N__1292),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1366),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1223));
    IO_PAD A_ibuf_0_iopad (
            .OE(N__2795),
            .DIN(N__2794),
            .DOUT(N__2793),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__2795),
            .PADOUT(N__2794),
            .PADIN(N__2793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_5_iopad (
            .OE(N__2786),
            .DIN(N__2785),
            .DOUT(N__2784),
            .PACKAGEPIN(B[5]));
    defparam B_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_5_preio (
            .PADOEN(N__2786),
            .PADOUT(N__2785),
            .PADIN(N__2784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_1_iopad (
            .OE(N__2777),
            .DIN(N__2776),
            .DOUT(N__2775),
            .PACKAGEPIN(alu_out[1]));
    defparam alu_out_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_1_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_1_preio (
            .PADOEN(N__2777),
            .PADOUT(N__2776),
            .PADIN(N__2775),
            .CLOCKENABLE(N__1297),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1225));
    IO_PAD s_ibuf_2_iopad (
            .OE(N__2768),
            .DIN(N__2767),
            .DOUT(N__2766),
            .PACKAGEPIN(s[2]));
    defparam s_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam s_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO s_ibuf_2_preio (
            .PADOEN(N__2768),
            .PADOUT(N__2767),
            .PADIN(N__2766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(s_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__2759),
            .DIN(N__2758),
            .DOUT(N__2757),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__2759),
            .PADOUT(N__2758),
            .PADIN(N__2757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_1_iopad (
            .OE(N__2750),
            .DIN(N__2749),
            .DOUT(N__2748),
            .PACKAGEPIN(B[1]));
    defparam B_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_1_preio (
            .PADOEN(N__2750),
            .PADOUT(N__2749),
            .PADIN(N__2748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD alu_out_obuf_5_iopad (
            .OE(N__2741),
            .DIN(N__2740),
            .DOUT(N__2739),
            .PACKAGEPIN(alu_out[5]));
    defparam alu_out_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam alu_out_obuf_5_preio.PIN_TYPE=6'b010101;
    PRE_IO alu_out_obuf_5_preio (
            .PADOEN(N__2741),
            .PADOUT(N__2740),
            .PADIN(N__2739),
            .CLOCKENABLE(N__1267),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1375),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1221));
    IO_PAD A_ibuf_1_iopad (
            .OE(N__2732),
            .DIN(N__2731),
            .DOUT(N__2730),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__2732),
            .PADOUT(N__2731),
            .PADIN(N__2730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_ibuf_4_iopad (
            .OE(N__2723),
            .DIN(N__2722),
            .DOUT(N__2721),
            .PACKAGEPIN(B[4]));
    defparam B_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam B_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO B_ibuf_4_preio (
            .PADOEN(N__2723),
            .PADOUT(N__2722),
            .PADIN(N__2721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(B_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s_ibuf_3_iopad (
            .OE(N__2714),
            .DIN(N__2713),
            .DOUT(N__2712),
            .PACKAGEPIN(s[3]));
    defparam s_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam s_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO s_ibuf_3_preio (
            .PADOEN(N__2714),
            .PADOUT(N__2713),
            .PADIN(N__2712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(s_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__601 (
            .O(N__2695),
            .I(alu_out_RNO_2Z0Z_6_cascade_));
    InMux I__600 (
            .O(N__2692),
            .I(N__2689));
    LocalMux I__599 (
            .O(N__2689),
            .I(alu_out_RNO_3Z0Z_6));
    InMux I__598 (
            .O(N__2686),
            .I(N__2683));
    LocalMux I__597 (
            .O(N__2683),
            .I(N__2680));
    Odrv4 I__596 (
            .O(N__2680),
            .I(N_148));
    CascadeMux I__595 (
            .O(N__2677),
            .I(N__2673));
    InMux I__594 (
            .O(N__2676),
            .I(N__2670));
    InMux I__593 (
            .O(N__2673),
            .I(N__2666));
    LocalMux I__592 (
            .O(N__2670),
            .I(N__2663));
    InMux I__591 (
            .O(N__2669),
            .I(N__2660));
    LocalMux I__590 (
            .O(N__2666),
            .I(N__2657));
    Span12Mux_s1_h I__589 (
            .O(N__2663),
            .I(N__2652));
    LocalMux I__588 (
            .O(N__2660),
            .I(N__2652));
    Odrv12 I__587 (
            .O(N__2657),
            .I(B_c_3));
    Odrv12 I__586 (
            .O(N__2652),
            .I(B_c_3));
    CascadeMux I__585 (
            .O(N__2647),
            .I(N__2644));
    InMux I__584 (
            .O(N__2644),
            .I(N__2637));
    InMux I__583 (
            .O(N__2643),
            .I(N__2637));
    CascadeMux I__582 (
            .O(N__2642),
            .I(N__2634));
    LocalMux I__581 (
            .O(N__2637),
            .I(N__2630));
    InMux I__580 (
            .O(N__2634),
            .I(N__2627));
    InMux I__579 (
            .O(N__2633),
            .I(N__2624));
    Span4Mux_v I__578 (
            .O(N__2630),
            .I(N__2619));
    LocalMux I__577 (
            .O(N__2627),
            .I(N__2619));
    LocalMux I__576 (
            .O(N__2624),
            .I(N__2616));
    Span4Mux_v I__575 (
            .O(N__2619),
            .I(N__2613));
    Span4Mux_v I__574 (
            .O(N__2616),
            .I(N__2610));
    Odrv4 I__573 (
            .O(N__2613),
            .I(A_c_3));
    Odrv4 I__572 (
            .O(N__2610),
            .I(A_c_3));
    CascadeMux I__571 (
            .O(N__2605),
            .I(N__2602));
    InMux I__570 (
            .O(N__2602),
            .I(N__2599));
    LocalMux I__569 (
            .O(N__2599),
            .I(N__2596));
    Odrv4 I__568 (
            .O(N__2596),
            .I(B_ibuf_RNI4CQF1Z0Z_3));
    CascadeMux I__567 (
            .O(N__2593),
            .I(N__2588));
    InMux I__566 (
            .O(N__2592),
            .I(N__2581));
    InMux I__565 (
            .O(N__2591),
            .I(N__2581));
    InMux I__564 (
            .O(N__2588),
            .I(N__2581));
    LocalMux I__563 (
            .O(N__2581),
            .I(N__2577));
    InMux I__562 (
            .O(N__2580),
            .I(N__2574));
    Odrv12 I__561 (
            .O(N__2577),
            .I(A_c_6));
    LocalMux I__560 (
            .O(N__2574),
            .I(A_c_6));
    InMux I__559 (
            .O(N__2569),
            .I(N__2564));
    InMux I__558 (
            .O(N__2568),
            .I(N__2559));
    InMux I__557 (
            .O(N__2567),
            .I(N__2559));
    LocalMux I__556 (
            .O(N__2564),
            .I(N__2556));
    LocalMux I__555 (
            .O(N__2559),
            .I(N__2553));
    Span4Mux_v I__554 (
            .O(N__2556),
            .I(N__2550));
    Span12Mux_s5_v I__553 (
            .O(N__2553),
            .I(N__2547));
    Odrv4 I__552 (
            .O(N__2550),
            .I(B_c_6));
    Odrv12 I__551 (
            .O(N__2547),
            .I(B_c_6));
    CascadeMux I__550 (
            .O(N__2542),
            .I(N__2539));
    InMux I__549 (
            .O(N__2539),
            .I(N__2536));
    LocalMux I__548 (
            .O(N__2536),
            .I(N__2533));
    Odrv4 I__547 (
            .O(N__2533),
            .I(B_ibuf_RNIAIQF1Z0Z_6));
    CascadeMux I__546 (
            .O(N__2530),
            .I(N__2525));
    InMux I__545 (
            .O(N__2529),
            .I(N__2520));
    InMux I__544 (
            .O(N__2528),
            .I(N__2520));
    InMux I__543 (
            .O(N__2525),
            .I(N__2517));
    LocalMux I__542 (
            .O(N__2520),
            .I(N__2514));
    LocalMux I__541 (
            .O(N__2517),
            .I(N__2510));
    Span4Mux_h I__540 (
            .O(N__2514),
            .I(N__2507));
    InMux I__539 (
            .O(N__2513),
            .I(N__2504));
    Span12Mux_s11_h I__538 (
            .O(N__2510),
            .I(N__2501));
    Span4Mux_v I__537 (
            .O(N__2507),
            .I(N__2498));
    LocalMux I__536 (
            .O(N__2504),
            .I(N__2495));
    Odrv12 I__535 (
            .O(N__2501),
            .I(A_c_7));
    Odrv4 I__534 (
            .O(N__2498),
            .I(A_c_7));
    Odrv12 I__533 (
            .O(N__2495),
            .I(A_c_7));
    InMux I__532 (
            .O(N__2488),
            .I(N__2469));
    InMux I__531 (
            .O(N__2487),
            .I(N__2469));
    InMux I__530 (
            .O(N__2486),
            .I(N__2469));
    InMux I__529 (
            .O(N__2485),
            .I(N__2469));
    InMux I__528 (
            .O(N__2484),
            .I(N__2466));
    InMux I__527 (
            .O(N__2483),
            .I(N__2459));
    InMux I__526 (
            .O(N__2482),
            .I(N__2459));
    InMux I__525 (
            .O(N__2481),
            .I(N__2459));
    InMux I__524 (
            .O(N__2480),
            .I(N__2452));
    InMux I__523 (
            .O(N__2479),
            .I(N__2452));
    InMux I__522 (
            .O(N__2478),
            .I(N__2452));
    LocalMux I__521 (
            .O(N__2469),
            .I(N__2446));
    LocalMux I__520 (
            .O(N__2466),
            .I(N__2446));
    LocalMux I__519 (
            .O(N__2459),
            .I(N__2441));
    LocalMux I__518 (
            .O(N__2452),
            .I(N__2441));
    CascadeMux I__517 (
            .O(N__2451),
            .I(N__2434));
    Span4Mux_v I__516 (
            .O(N__2446),
            .I(N__2428));
    Span4Mux_v I__515 (
            .O(N__2441),
            .I(N__2425));
    InMux I__514 (
            .O(N__2440),
            .I(N__2418));
    InMux I__513 (
            .O(N__2439),
            .I(N__2418));
    InMux I__512 (
            .O(N__2438),
            .I(N__2418));
    InMux I__511 (
            .O(N__2437),
            .I(N__2411));
    InMux I__510 (
            .O(N__2434),
            .I(N__2411));
    InMux I__509 (
            .O(N__2433),
            .I(N__2411));
    InMux I__508 (
            .O(N__2432),
            .I(N__2406));
    InMux I__507 (
            .O(N__2431),
            .I(N__2406));
    Sp12to4 I__506 (
            .O(N__2428),
            .I(N__2399));
    Sp12to4 I__505 (
            .O(N__2425),
            .I(N__2399));
    LocalMux I__504 (
            .O(N__2418),
            .I(N__2399));
    LocalMux I__503 (
            .O(N__2411),
            .I(s_c_1));
    LocalMux I__502 (
            .O(N__2406),
            .I(s_c_1));
    Odrv12 I__501 (
            .O(N__2399),
            .I(s_c_1));
    CascadeMux I__500 (
            .O(N__2392),
            .I(N__2386));
    CascadeMux I__499 (
            .O(N__2391),
            .I(N__2383));
    CascadeMux I__498 (
            .O(N__2390),
            .I(N__2368));
    InMux I__497 (
            .O(N__2389),
            .I(N__2352));
    InMux I__496 (
            .O(N__2386),
            .I(N__2352));
    InMux I__495 (
            .O(N__2383),
            .I(N__2352));
    InMux I__494 (
            .O(N__2382),
            .I(N__2352));
    InMux I__493 (
            .O(N__2381),
            .I(N__2347));
    InMux I__492 (
            .O(N__2380),
            .I(N__2347));
    InMux I__491 (
            .O(N__2379),
            .I(N__2338));
    InMux I__490 (
            .O(N__2378),
            .I(N__2338));
    InMux I__489 (
            .O(N__2377),
            .I(N__2338));
    InMux I__488 (
            .O(N__2376),
            .I(N__2338));
    InMux I__487 (
            .O(N__2375),
            .I(N__2327));
    InMux I__486 (
            .O(N__2374),
            .I(N__2327));
    InMux I__485 (
            .O(N__2373),
            .I(N__2327));
    InMux I__484 (
            .O(N__2372),
            .I(N__2327));
    InMux I__483 (
            .O(N__2371),
            .I(N__2327));
    InMux I__482 (
            .O(N__2368),
            .I(N__2318));
    InMux I__481 (
            .O(N__2367),
            .I(N__2318));
    InMux I__480 (
            .O(N__2366),
            .I(N__2318));
    InMux I__479 (
            .O(N__2365),
            .I(N__2318));
    InMux I__478 (
            .O(N__2364),
            .I(N__2309));
    InMux I__477 (
            .O(N__2363),
            .I(N__2309));
    InMux I__476 (
            .O(N__2362),
            .I(N__2309));
    InMux I__475 (
            .O(N__2361),
            .I(N__2309));
    LocalMux I__474 (
            .O(N__2352),
            .I(N__2304));
    LocalMux I__473 (
            .O(N__2347),
            .I(N__2297));
    LocalMux I__472 (
            .O(N__2338),
            .I(N__2297));
    LocalMux I__471 (
            .O(N__2327),
            .I(N__2297));
    LocalMux I__470 (
            .O(N__2318),
            .I(N__2292));
    LocalMux I__469 (
            .O(N__2309),
            .I(N__2292));
    CascadeMux I__468 (
            .O(N__2308),
            .I(N__2280));
    CascadeMux I__467 (
            .O(N__2307),
            .I(N__2275));
    Span4Mux_v I__466 (
            .O(N__2304),
            .I(N__2268));
    Span4Mux_v I__465 (
            .O(N__2297),
            .I(N__2268));
    Span4Mux_v I__464 (
            .O(N__2292),
            .I(N__2268));
    InMux I__463 (
            .O(N__2291),
            .I(N__2259));
    InMux I__462 (
            .O(N__2290),
            .I(N__2259));
    InMux I__461 (
            .O(N__2289),
            .I(N__2259));
    InMux I__460 (
            .O(N__2288),
            .I(N__2259));
    InMux I__459 (
            .O(N__2287),
            .I(N__2246));
    InMux I__458 (
            .O(N__2286),
            .I(N__2246));
    InMux I__457 (
            .O(N__2285),
            .I(N__2246));
    InMux I__456 (
            .O(N__2284),
            .I(N__2246));
    InMux I__455 (
            .O(N__2283),
            .I(N__2246));
    InMux I__454 (
            .O(N__2280),
            .I(N__2246));
    InMux I__453 (
            .O(N__2279),
            .I(N__2239));
    InMux I__452 (
            .O(N__2278),
            .I(N__2239));
    InMux I__451 (
            .O(N__2275),
            .I(N__2239));
    Odrv4 I__450 (
            .O(N__2268),
            .I(s_c_0));
    LocalMux I__449 (
            .O(N__2259),
            .I(s_c_0));
    LocalMux I__448 (
            .O(N__2246),
            .I(s_c_0));
    LocalMux I__447 (
            .O(N__2239),
            .I(s_c_0));
    InMux I__446 (
            .O(N__2230),
            .I(N__2225));
    InMux I__445 (
            .O(N__2229),
            .I(N__2222));
    InMux I__444 (
            .O(N__2228),
            .I(N__2219));
    LocalMux I__443 (
            .O(N__2225),
            .I(N__2216));
    LocalMux I__442 (
            .O(N__2222),
            .I(N__2211));
    LocalMux I__441 (
            .O(N__2219),
            .I(N__2211));
    Span4Mux_v I__440 (
            .O(N__2216),
            .I(N__2208));
    Odrv12 I__439 (
            .O(N__2211),
            .I(B_c_7));
    Odrv4 I__438 (
            .O(N__2208),
            .I(B_c_7));
    InMux I__437 (
            .O(N__2203),
            .I(N__2192));
    InMux I__436 (
            .O(N__2202),
            .I(N__2192));
    InMux I__435 (
            .O(N__2201),
            .I(N__2189));
    InMux I__434 (
            .O(N__2200),
            .I(N__2184));
    InMux I__433 (
            .O(N__2199),
            .I(N__2184));
    InMux I__432 (
            .O(N__2198),
            .I(N__2179));
    InMux I__431 (
            .O(N__2197),
            .I(N__2179));
    LocalMux I__430 (
            .O(N__2192),
            .I(N__2174));
    LocalMux I__429 (
            .O(N__2189),
            .I(N__2174));
    LocalMux I__428 (
            .O(N__2184),
            .I(N__2169));
    LocalMux I__427 (
            .O(N__2179),
            .I(N__2169));
    Span4Mux_v I__426 (
            .O(N__2174),
            .I(N__2162));
    Span4Mux_v I__425 (
            .O(N__2169),
            .I(N__2159));
    InMux I__424 (
            .O(N__2168),
            .I(N__2150));
    InMux I__423 (
            .O(N__2167),
            .I(N__2150));
    InMux I__422 (
            .O(N__2166),
            .I(N__2150));
    InMux I__421 (
            .O(N__2165),
            .I(N__2150));
    Odrv4 I__420 (
            .O(N__2162),
            .I(s_c_2));
    Odrv4 I__419 (
            .O(N__2159),
            .I(s_c_2));
    LocalMux I__418 (
            .O(N__2150),
            .I(s_c_2));
    InMux I__417 (
            .O(N__2143),
            .I(N__2140));
    LocalMux I__416 (
            .O(N__2140),
            .I(alu_out_RNO_5Z0Z_7));
    CascadeMux I__415 (
            .O(N__2137),
            .I(alu_out_RNO_4Z0Z_7_cascade_));
    InMux I__414 (
            .O(N__2134),
            .I(N__2131));
    LocalMux I__413 (
            .O(N__2131),
            .I(N_149));
    InMux I__412 (
            .O(N__2128),
            .I(N__2125));
    LocalMux I__411 (
            .O(N__2125),
            .I(alu_out_RNO_3Z0Z_7));
    InMux I__410 (
            .O(N__2122),
            .I(N__2119));
    LocalMux I__409 (
            .O(N__2119),
            .I(N_91));
    InMux I__408 (
            .O(N__2116),
            .I(N__2113));
    LocalMux I__407 (
            .O(N__2113),
            .I(N__2110));
    Odrv4 I__406 (
            .O(N__2110),
            .I(B_ibuf_RNII15C1Z0Z_2));
    CascadeMux I__405 (
            .O(N__2107),
            .I(N__2103));
    InMux I__404 (
            .O(N__2106),
            .I(N__2098));
    InMux I__403 (
            .O(N__2103),
            .I(N__2098));
    LocalMux I__402 (
            .O(N__2098),
            .I(N__2094));
    InMux I__401 (
            .O(N__2097),
            .I(N__2091));
    Span4Mux_v I__400 (
            .O(N__2094),
            .I(N__2086));
    LocalMux I__399 (
            .O(N__2091),
            .I(N__2086));
    Span4Mux_v I__398 (
            .O(N__2086),
            .I(N__2083));
    Odrv4 I__397 (
            .O(N__2083),
            .I(B_c_2));
    InMux I__396 (
            .O(N__2080),
            .I(N__2077));
    LocalMux I__395 (
            .O(N__2077),
            .I(N_86));
    InMux I__394 (
            .O(N__2074),
            .I(N__2071));
    LocalMux I__393 (
            .O(N__2071),
            .I(N__2067));
    CascadeMux I__392 (
            .O(N__2070),
            .I(N__2064));
    Span4Mux_v I__391 (
            .O(N__2067),
            .I(N__2060));
    InMux I__390 (
            .O(N__2064),
            .I(N__2055));
    InMux I__389 (
            .O(N__2063),
            .I(N__2055));
    Odrv4 I__388 (
            .O(N__2060),
            .I(B_c_5));
    LocalMux I__387 (
            .O(N__2055),
            .I(B_c_5));
    CascadeMux I__386 (
            .O(N__2050),
            .I(N_89_cascade_));
    InMux I__385 (
            .O(N__2047),
            .I(N__2044));
    LocalMux I__384 (
            .O(N__2044),
            .I(B_ibuf_RNIL45C1Z0Z_5));
    InMux I__383 (
            .O(N__2041),
            .I(N__2035));
    InMux I__382 (
            .O(N__2040),
            .I(N__2027));
    InMux I__381 (
            .O(N__2039),
            .I(N__2027));
    CascadeMux I__380 (
            .O(N__2038),
            .I(N__2022));
    LocalMux I__379 (
            .O(N__2035),
            .I(N__2016));
    InMux I__378 (
            .O(N__2034),
            .I(N__2009));
    InMux I__377 (
            .O(N__2033),
            .I(N__2009));
    InMux I__376 (
            .O(N__2032),
            .I(N__2009));
    LocalMux I__375 (
            .O(N__2027),
            .I(N__2006));
    InMux I__374 (
            .O(N__2026),
            .I(N__2001));
    InMux I__373 (
            .O(N__2025),
            .I(N__2001));
    InMux I__372 (
            .O(N__2022),
            .I(N__1994));
    InMux I__371 (
            .O(N__2021),
            .I(N__1994));
    InMux I__370 (
            .O(N__2020),
            .I(N__1994));
    InMux I__369 (
            .O(N__2019),
            .I(N__1991));
    Odrv4 I__368 (
            .O(N__2016),
            .I(s_c_i_1));
    LocalMux I__367 (
            .O(N__2009),
            .I(s_c_i_1));
    Odrv4 I__366 (
            .O(N__2006),
            .I(s_c_i_1));
    LocalMux I__365 (
            .O(N__2001),
            .I(s_c_i_1));
    LocalMux I__364 (
            .O(N__1994),
            .I(s_c_i_1));
    LocalMux I__363 (
            .O(N__1991),
            .I(s_c_i_1));
    CascadeMux I__362 (
            .O(N__1978),
            .I(N__1975));
    InMux I__361 (
            .O(N__1975),
            .I(N__1971));
    InMux I__360 (
            .O(N__1974),
            .I(N__1968));
    LocalMux I__359 (
            .O(N__1971),
            .I(N__1965));
    LocalMux I__358 (
            .O(N__1968),
            .I(N__1962));
    Span4Mux_v I__357 (
            .O(N__1965),
            .I(N__1957));
    Span4Mux_v I__356 (
            .O(N__1962),
            .I(N__1954));
    InMux I__355 (
            .O(N__1961),
            .I(N__1949));
    InMux I__354 (
            .O(N__1960),
            .I(N__1949));
    Odrv4 I__353 (
            .O(N__1957),
            .I(A_c_0));
    Odrv4 I__352 (
            .O(N__1954),
            .I(A_c_0));
    LocalMux I__351 (
            .O(N__1949),
            .I(A_c_0));
    InMux I__350 (
            .O(N__1942),
            .I(N__1939));
    LocalMux I__349 (
            .O(N__1939),
            .I(N__1935));
    CascadeMux I__348 (
            .O(N__1938),
            .I(N__1930));
    Span4Mux_v I__347 (
            .O(N__1935),
            .I(N__1927));
    InMux I__346 (
            .O(N__1934),
            .I(N__1924));
    InMux I__345 (
            .O(N__1933),
            .I(N__1919));
    InMux I__344 (
            .O(N__1930),
            .I(N__1919));
    Odrv4 I__343 (
            .O(N__1927),
            .I(A_c_5));
    LocalMux I__342 (
            .O(N__1924),
            .I(A_c_5));
    LocalMux I__341 (
            .O(N__1919),
            .I(A_c_5));
    InMux I__340 (
            .O(N__1912),
            .I(N__1909));
    LocalMux I__339 (
            .O(N__1909),
            .I(B_ibuf_RNIH05C1Z0Z_1));
    CascadeMux I__338 (
            .O(N__1906),
            .I(N__1903));
    InMux I__337 (
            .O(N__1903),
            .I(N__1900));
    LocalMux I__336 (
            .O(N__1900),
            .I(B_ibuf_RNI08QF1Z0Z_1));
    InMux I__335 (
            .O(N__1897),
            .I(N__1894));
    LocalMux I__334 (
            .O(N__1894),
            .I(N__1891));
    Odrv4 I__333 (
            .O(N__1891),
            .I(alu_out_RNO_1Z0Z_1));
    InMux I__332 (
            .O(N__1888),
            .I(un1_A_1_cry_0));
    CascadeMux I__331 (
            .O(N__1885),
            .I(N__1882));
    InMux I__330 (
            .O(N__1882),
            .I(N__1879));
    LocalMux I__329 (
            .O(N__1879),
            .I(B_ibuf_RNI2AQF1Z0Z_2));
    InMux I__328 (
            .O(N__1876),
            .I(N__1873));
    LocalMux I__327 (
            .O(N__1873),
            .I(alu_out_RNO_1Z0Z_2));
    InMux I__326 (
            .O(N__1870),
            .I(un1_A_1_cry_1));
    InMux I__325 (
            .O(N__1867),
            .I(N__1864));
    LocalMux I__324 (
            .O(N__1864),
            .I(B_ibuf_RNIJ25C1Z0Z_3));
    InMux I__323 (
            .O(N__1861),
            .I(N__1858));
    LocalMux I__322 (
            .O(N__1858),
            .I(alu_out_RNO_1Z0Z_3));
    InMux I__321 (
            .O(N__1855),
            .I(un1_A_1_cry_2));
    InMux I__320 (
            .O(N__1852),
            .I(N__1849));
    LocalMux I__319 (
            .O(N__1849),
            .I(B_ibuf_RNIK35C1Z0Z_4));
    CascadeMux I__318 (
            .O(N__1846),
            .I(N__1843));
    InMux I__317 (
            .O(N__1843),
            .I(N__1840));
    LocalMux I__316 (
            .O(N__1840),
            .I(B_ibuf_RNI6EQF1Z0Z_4));
    InMux I__315 (
            .O(N__1837),
            .I(N__1834));
    LocalMux I__314 (
            .O(N__1834),
            .I(alu_out_RNO_1Z0Z_4));
    InMux I__313 (
            .O(N__1831),
            .I(un1_A_1_cry_3));
    CascadeMux I__312 (
            .O(N__1828),
            .I(N__1825));
    InMux I__311 (
            .O(N__1825),
            .I(N__1822));
    LocalMux I__310 (
            .O(N__1822),
            .I(N__1819));
    Odrv4 I__309 (
            .O(N__1819),
            .I(B_ibuf_RNI8GQF1Z0Z_5));
    InMux I__308 (
            .O(N__1816),
            .I(N__1813));
    LocalMux I__307 (
            .O(N__1813),
            .I(alu_out_RNO_1Z0Z_5));
    InMux I__306 (
            .O(N__1810),
            .I(un1_A_1_cry_4));
    InMux I__305 (
            .O(N__1807),
            .I(N__1804));
    LocalMux I__304 (
            .O(N__1804),
            .I(N__1801));
    Odrv4 I__303 (
            .O(N__1801),
            .I(B_ibuf_RNIM55C1Z0Z_6));
    InMux I__302 (
            .O(N__1798),
            .I(N__1795));
    LocalMux I__301 (
            .O(N__1795),
            .I(alu_out_RNO_1Z0Z_6));
    InMux I__300 (
            .O(N__1792),
            .I(un1_A_1_cry_5));
    CascadeMux I__299 (
            .O(N__1789),
            .I(N__1786));
    InMux I__298 (
            .O(N__1786),
            .I(N__1783));
    LocalMux I__297 (
            .O(N__1783),
            .I(N__1774));
    InMux I__296 (
            .O(N__1782),
            .I(N__1769));
    InMux I__295 (
            .O(N__1781),
            .I(N__1769));
    InMux I__294 (
            .O(N__1780),
            .I(N__1760));
    InMux I__293 (
            .O(N__1779),
            .I(N__1760));
    InMux I__292 (
            .O(N__1778),
            .I(N__1760));
    InMux I__291 (
            .O(N__1777),
            .I(N__1760));
    Span4Mux_v I__290 (
            .O(N__1774),
            .I(N__1755));
    LocalMux I__289 (
            .O(N__1769),
            .I(N__1755));
    LocalMux I__288 (
            .O(N__1760),
            .I(N__1752));
    Span4Mux_v I__287 (
            .O(N__1755),
            .I(N__1745));
    Span4Mux_v I__286 (
            .O(N__1752),
            .I(N__1742));
    InMux I__285 (
            .O(N__1751),
            .I(N__1739));
    InMux I__284 (
            .O(N__1750),
            .I(N__1732));
    InMux I__283 (
            .O(N__1749),
            .I(N__1732));
    InMux I__282 (
            .O(N__1748),
            .I(N__1732));
    Odrv4 I__281 (
            .O(N__1745),
            .I(s_c_3));
    Odrv4 I__280 (
            .O(N__1742),
            .I(s_c_3));
    LocalMux I__279 (
            .O(N__1739),
            .I(s_c_3));
    LocalMux I__278 (
            .O(N__1732),
            .I(s_c_3));
    InMux I__277 (
            .O(N__1723),
            .I(bfn_2_11_0_));
    IoInMux I__276 (
            .O(N__1720),
            .I(N__1717));
    LocalMux I__275 (
            .O(N__1717),
            .I(N__1714));
    IoSpan4Mux I__274 (
            .O(N__1714),
            .I(N__1711));
    Span4Mux_s1_h I__273 (
            .O(N__1711),
            .I(N__1708));
    Span4Mux_h I__272 (
            .O(N__1708),
            .I(N__1705));
    Odrv4 I__271 (
            .O(N__1705),
            .I(alu_out_13_7));
    InMux I__270 (
            .O(N__1702),
            .I(N__1699));
    LocalMux I__269 (
            .O(N__1699),
            .I(un1_A_1_axb_7));
    CascadeMux I__268 (
            .O(N__1696),
            .I(alu_out_RNO_2Z0Z_3_cascade_));
    InMux I__267 (
            .O(N__1693),
            .I(N__1690));
    LocalMux I__266 (
            .O(N__1690),
            .I(alu_out_RNO_3Z0Z_3));
    CascadeMux I__265 (
            .O(N__1687),
            .I(N_145_cascade_));
    IoInMux I__264 (
            .O(N__1684),
            .I(N__1681));
    LocalMux I__263 (
            .O(N__1681),
            .I(N__1678));
    Span4Mux_s2_h I__262 (
            .O(N__1678),
            .I(N__1675));
    Odrv4 I__261 (
            .O(N__1675),
            .I(alu_out_13_3));
    CascadeMux I__260 (
            .O(N__1672),
            .I(N__1669));
    InMux I__259 (
            .O(N__1669),
            .I(N__1661));
    InMux I__258 (
            .O(N__1668),
            .I(N__1661));
    InMux I__257 (
            .O(N__1667),
            .I(N__1656));
    InMux I__256 (
            .O(N__1666),
            .I(N__1656));
    LocalMux I__255 (
            .O(N__1661),
            .I(N__1651));
    LocalMux I__254 (
            .O(N__1656),
            .I(N__1651));
    Span4Mux_v I__253 (
            .O(N__1651),
            .I(N__1648));
    Span4Mux_v I__252 (
            .O(N__1648),
            .I(N__1645));
    Odrv4 I__251 (
            .O(N__1645),
            .I(A_c_2));
    InMux I__250 (
            .O(N__1642),
            .I(N__1634));
    InMux I__249 (
            .O(N__1641),
            .I(N__1634));
    InMux I__248 (
            .O(N__1640),
            .I(N__1631));
    InMux I__247 (
            .O(N__1639),
            .I(N__1628));
    LocalMux I__246 (
            .O(N__1634),
            .I(N__1621));
    LocalMux I__245 (
            .O(N__1631),
            .I(N__1621));
    LocalMux I__244 (
            .O(N__1628),
            .I(N__1621));
    Span4Mux_v I__243 (
            .O(N__1621),
            .I(N__1618));
    Span4Mux_v I__242 (
            .O(N__1618),
            .I(N__1615));
    Odrv4 I__241 (
            .O(N__1615),
            .I(A_c_1));
    CascadeMux I__240 (
            .O(N__1612),
            .I(alu_out_RNO_3Z0Z_2_cascade_));
    InMux I__239 (
            .O(N__1609),
            .I(N__1606));
    LocalMux I__238 (
            .O(N__1606),
            .I(alu_out_RNO_2Z0Z_2));
    CascadeMux I__237 (
            .O(N__1603),
            .I(N_144_cascade_));
    IoInMux I__236 (
            .O(N__1600),
            .I(N__1597));
    LocalMux I__235 (
            .O(N__1597),
            .I(N__1594));
    Span12Mux_s1_h I__234 (
            .O(N__1594),
            .I(N__1591));
    Odrv12 I__233 (
            .O(N__1591),
            .I(alu_out_13_2));
    CascadeMux I__232 (
            .O(N__1588),
            .I(N__1585));
    InMux I__231 (
            .O(N__1585),
            .I(N__1581));
    InMux I__230 (
            .O(N__1584),
            .I(N__1578));
    LocalMux I__229 (
            .O(N__1581),
            .I(s_ibuf_RNI1HJVZ0Z_0));
    LocalMux I__228 (
            .O(N__1578),
            .I(s_ibuf_RNI1HJVZ0Z_0));
    InMux I__227 (
            .O(N__1573),
            .I(N__1570));
    LocalMux I__226 (
            .O(N__1570),
            .I(un1_A_1));
    CascadeMux I__225 (
            .O(N__1567),
            .I(N__1564));
    InMux I__224 (
            .O(N__1564),
            .I(N__1561));
    LocalMux I__223 (
            .O(N__1561),
            .I(B_ibuf_RNIE5VR2Z0Z_0));
    InMux I__222 (
            .O(N__1558),
            .I(N__1555));
    LocalMux I__221 (
            .O(N__1555),
            .I(alu_out_RNO_1Z0Z_0));
    InMux I__220 (
            .O(N__1552),
            .I(un1_A_1_cry_0_c_THRU_CO));
    CascadeMux I__219 (
            .O(N__1549),
            .I(N_85_cascade_));
    InMux I__218 (
            .O(N__1546),
            .I(N__1540));
    InMux I__217 (
            .O(N__1545),
            .I(N__1540));
    LocalMux I__216 (
            .O(N__1540),
            .I(N__1536));
    CascadeMux I__215 (
            .O(N__1539),
            .I(N__1533));
    Span4Mux_v I__214 (
            .O(N__1536),
            .I(N__1530));
    InMux I__213 (
            .O(N__1533),
            .I(N__1527));
    Odrv4 I__212 (
            .O(N__1530),
            .I(B_c_4));
    LocalMux I__211 (
            .O(N__1527),
            .I(B_c_4));
    InMux I__210 (
            .O(N__1522),
            .I(N__1519));
    LocalMux I__209 (
            .O(N__1519),
            .I(alu_out_RNO_3Z0Z_4));
    CascadeMux I__208 (
            .O(N__1516),
            .I(alu_out_RNO_2Z0Z_4_cascade_));
    InMux I__207 (
            .O(N__1513),
            .I(N__1510));
    LocalMux I__206 (
            .O(N__1510),
            .I(N__1507));
    Odrv4 I__205 (
            .O(N__1507),
            .I(N_146));
    InMux I__204 (
            .O(N__1504),
            .I(N__1500));
    InMux I__203 (
            .O(N__1503),
            .I(N__1497));
    LocalMux I__202 (
            .O(N__1500),
            .I(N__1492));
    LocalMux I__201 (
            .O(N__1497),
            .I(N__1489));
    InMux I__200 (
            .O(N__1496),
            .I(N__1484));
    InMux I__199 (
            .O(N__1495),
            .I(N__1484));
    Span4Mux_v I__198 (
            .O(N__1492),
            .I(N__1477));
    Span4Mux_h I__197 (
            .O(N__1489),
            .I(N__1477));
    LocalMux I__196 (
            .O(N__1484),
            .I(N__1477));
    Span4Mux_v I__195 (
            .O(N__1477),
            .I(N__1474));
    Odrv4 I__194 (
            .O(N__1474),
            .I(A_c_4));
    CascadeMux I__193 (
            .O(N__1471),
            .I(alu_out_RNO_2Z0Z_5_cascade_));
    InMux I__192 (
            .O(N__1468),
            .I(N__1465));
    LocalMux I__191 (
            .O(N__1465),
            .I(alu_out_RNO_3Z0Z_5));
    InMux I__190 (
            .O(N__1462),
            .I(N__1459));
    LocalMux I__189 (
            .O(N__1459),
            .I(N__1456));
    Odrv12 I__188 (
            .O(N__1456),
            .I(N_147));
    CascadeMux I__187 (
            .O(N__1453),
            .I(s_c_i_1_cascade_));
    InMux I__186 (
            .O(N__1450),
            .I(N__1447));
    LocalMux I__185 (
            .O(N__1447),
            .I(N_88));
    CascadeMux I__184 (
            .O(N__1444),
            .I(un1_A_1_cascade_));
    CascadeMux I__183 (
            .O(N__1441),
            .I(N__1437));
    CascadeMux I__182 (
            .O(N__1440),
            .I(N__1434));
    InMux I__181 (
            .O(N__1437),
            .I(N__1426));
    InMux I__180 (
            .O(N__1434),
            .I(N__1426));
    InMux I__179 (
            .O(N__1433),
            .I(N__1426));
    LocalMux I__178 (
            .O(N__1426),
            .I(N__1423));
    Odrv12 I__177 (
            .O(N__1423),
            .I(B_c_0));
    CascadeMux I__176 (
            .O(N__1420),
            .I(alu_out_RNO_2Z0Z_0_cascade_));
    InMux I__175 (
            .O(N__1417),
            .I(N__1414));
    LocalMux I__174 (
            .O(N__1414),
            .I(N_142));
    InMux I__173 (
            .O(N__1411),
            .I(N__1408));
    LocalMux I__172 (
            .O(N__1408),
            .I(alu_out_RNO_3Z0Z_0));
    InMux I__171 (
            .O(N__1405),
            .I(N__1398));
    InMux I__170 (
            .O(N__1404),
            .I(N__1398));
    CascadeMux I__169 (
            .O(N__1403),
            .I(N__1395));
    LocalMux I__168 (
            .O(N__1398),
            .I(N__1392));
    InMux I__167 (
            .O(N__1395),
            .I(N__1389));
    Span4Mux_v I__166 (
            .O(N__1392),
            .I(N__1384));
    LocalMux I__165 (
            .O(N__1389),
            .I(N__1384));
    Span4Mux_v I__164 (
            .O(N__1384),
            .I(N__1381));
    Span4Mux_v I__163 (
            .O(N__1381),
            .I(N__1378));
    Odrv4 I__162 (
            .O(N__1378),
            .I(B_c_1));
    IoInMux I__161 (
            .O(N__1375),
            .I(N__1372));
    LocalMux I__160 (
            .O(N__1372),
            .I(alu_out_13_5));
    CascadeMux I__159 (
            .O(N__1369),
            .I(N_87_cascade_));
    IoInMux I__158 (
            .O(N__1366),
            .I(N__1363));
    LocalMux I__157 (
            .O(N__1363),
            .I(N__1360));
    IoSpan4Mux I__156 (
            .O(N__1360),
            .I(N__1357));
    Span4Mux_s0_h I__155 (
            .O(N__1357),
            .I(N__1354));
    Odrv4 I__154 (
            .O(N__1354),
            .I(alu_out_13_4));
    IoInMux I__153 (
            .O(N__1351),
            .I(N__1348));
    LocalMux I__152 (
            .O(N__1348),
            .I(N__1345));
    IoSpan4Mux I__151 (
            .O(N__1345),
            .I(N__1342));
    Span4Mux_s0_h I__150 (
            .O(N__1342),
            .I(N__1339));
    Odrv4 I__149 (
            .O(N__1339),
            .I(alu_out_13_0));
    IoInMux I__148 (
            .O(N__1336),
            .I(N__1333));
    LocalMux I__147 (
            .O(N__1333),
            .I(N__1330));
    Span4Mux_s0_h I__146 (
            .O(N__1330),
            .I(N__1327));
    Span4Mux_v I__145 (
            .O(N__1327),
            .I(N__1324));
    Odrv4 I__144 (
            .O(N__1324),
            .I(alu_out_13_6));
    CascadeMux I__143 (
            .O(N__1321),
            .I(N_143_cascade_));
    IoInMux I__142 (
            .O(N__1318),
            .I(N__1315));
    LocalMux I__141 (
            .O(N__1315),
            .I(N__1312));
    Span4Mux_s0_h I__140 (
            .O(N__1312),
            .I(N__1309));
    Span4Mux_v I__139 (
            .O(N__1309),
            .I(N__1306));
    Odrv4 I__138 (
            .O(N__1306),
            .I(alu_out_13_1));
    CascadeMux I__137 (
            .O(N__1303),
            .I(alu_out38_cascade_));
    CascadeMux I__136 (
            .O(N__1300),
            .I(un1_alu_out43_1_3_cascade_));
    CEMux I__135 (
            .O(N__1297),
            .I(N__1293));
    CEMux I__134 (
            .O(N__1296),
            .I(N__1288));
    LocalMux I__133 (
            .O(N__1293),
            .I(N__1285));
    CEMux I__132 (
            .O(N__1292),
            .I(N__1282));
    CEMux I__131 (
            .O(N__1291),
            .I(N__1279));
    LocalMux I__130 (
            .O(N__1288),
            .I(N__1276));
    IoSpan4Mux I__129 (
            .O(N__1285),
            .I(N__1271));
    LocalMux I__128 (
            .O(N__1282),
            .I(N__1271));
    LocalMux I__127 (
            .O(N__1279),
            .I(N__1268));
    Span4Mux_s1_h I__126 (
            .O(N__1276),
            .I(N__1264));
    IoSpan4Mux I__125 (
            .O(N__1271),
            .I(N__1261));
    Span4Mux_s0_h I__124 (
            .O(N__1268),
            .I(N__1258));
    CEMux I__123 (
            .O(N__1267),
            .I(N__1255));
    Odrv4 I__122 (
            .O(N__1264),
            .I(un1_alu_out43_1_i));
    Odrv4 I__121 (
            .O(N__1261),
            .I(un1_alu_out43_1_i));
    Odrv4 I__120 (
            .O(N__1258),
            .I(un1_alu_out43_1_i));
    LocalMux I__119 (
            .O(N__1255),
            .I(un1_alu_out43_1_i));
    InMux I__118 (
            .O(N__1246),
            .I(N__1243));
    LocalMux I__117 (
            .O(N__1243),
            .I(un1_alu_out43_1_2));
    InMux I__116 (
            .O(N__1240),
            .I(N__1237));
    LocalMux I__115 (
            .O(N__1237),
            .I(alu_out40_0));
    CascadeMux I__114 (
            .O(N__1234),
            .I(N_90_cascade_));
    InMux I__113 (
            .O(N__1231),
            .I(N__1228));
    LocalMux I__112 (
            .O(N__1228),
            .I(alu_out_RNO_3Z0Z_1));
    ClkMux I__111 (
            .O(N__1225),
            .I(N__1210));
    ClkMux I__110 (
            .O(N__1224),
            .I(N__1210));
    ClkMux I__109 (
            .O(N__1223),
            .I(N__1210));
    ClkMux I__108 (
            .O(N__1222),
            .I(N__1210));
    ClkMux I__107 (
            .O(N__1221),
            .I(N__1210));
    GlobalMux I__106 (
            .O(N__1210),
            .I(N__1207));
    gio2CtrlBuf I__105 (
            .O(N__1207),
            .I(clk_c_g));
    CascadeMux I__104 (
            .O(N__1204),
            .I(alu_out_RNO_2Z0Z_1_cascade_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(un1_A_1_cry_6),
            .carryinitout(bfn_2_11_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam alu_out_RNO_2_1_LC_1_8_0.C_ON=1'b0;
    defparam alu_out_RNO_2_1_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_1_LC_1_8_0.LUT_INIT=16'b0101111001101000;
    LogicCell40 alu_out_RNO_2_1_LC_1_8_0 (
            .in0(N__2365),
            .in1(N__2433),
            .in2(N__1403),
            .in3(N__1639),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_1_LC_1_8_1.C_ON=1'b0;
    defparam alu_out_RNO_0_1_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_1_LC_1_8_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 alu_out_RNO_0_1_LC_1_8_1 (
            .in0(N__2165),
            .in1(_gnd_net_),
            .in2(N__1204),
            .in3(N__1231),
            .lcout(),
            .ltout(N_143_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_LC_1_8_2.C_ON=1'b0;
    defparam alu_out_RNO_1_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_LC_1_8_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 alu_out_RNO_1_LC_1_8_2 (
            .in0(N__1777),
            .in1(_gnd_net_),
            .in2(N__1321),
            .in3(N__1897),
            .lcout(alu_out_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNI667V1_0_2_LC_1_8_3.C_ON=1'b0;
    defparam s_ibuf_RNI667V1_0_2_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNI667V1_0_2_LC_1_8_3.LUT_INIT=16'b0000000001000000;
    LogicCell40 s_ibuf_RNI667V1_0_2_LC_1_8_3 (
            .in0(N__2166),
            .in1(N__1779),
            .in2(N__2451),
            .in3(N__2367),
            .lcout(),
            .ltout(alu_out38_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNID58E4_2_LC_1_8_4.C_ON=1'b0;
    defparam s_ibuf_RNID58E4_2_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNID58E4_2_LC_1_8_4.LUT_INIT=16'b0000010100000011;
    LogicCell40 s_ibuf_RNID58E4_2_LC_1_8_4 (
            .in0(N__1240),
            .in1(N__2040),
            .in2(N__1303),
            .in3(N__2168),
            .lcout(),
            .ltout(un1_alu_out43_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNIJBFD6_2_LC_1_8_5.C_ON=1'b0;
    defparam s_ibuf_RNIJBFD6_2_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNIJBFD6_2_LC_1_8_5.LUT_INIT=16'b0000111111111111;
    LogicCell40 s_ibuf_RNIJBFD6_2_LC_1_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1300),
            .in3(N__1246),
            .lcout(un1_alu_out43_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNI667V1_2_LC_1_8_6.C_ON=1'b0;
    defparam s_ibuf_RNI667V1_2_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNI667V1_2_LC_1_8_6.LUT_INIT=16'b0100011101110111;
    LogicCell40 s_ibuf_RNI667V1_2_LC_1_8_6 (
            .in0(N__1780),
            .in1(N__2167),
            .in2(N__2390),
            .in3(N__2437),
            .lcout(un1_alu_out43_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNI4CDF1_3_LC_1_8_7.C_ON=1'b0;
    defparam s_ibuf_RNI4CDF1_3_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNI4CDF1_3_LC_1_8_7.LUT_INIT=16'b0000000010001000;
    LogicCell40 s_ibuf_RNI4CDF1_3_LC_1_8_7 (
            .in0(N__2039),
            .in1(N__1778),
            .in2(_gnd_net_),
            .in3(N__2366),
            .lcout(alu_out40_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNILCBS_6_LC_1_9_0.C_ON=1'b0;
    defparam B_ibuf_RNILCBS_6_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNILCBS_6_LC_1_9_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 B_ibuf_RNILCBS_6_LC_1_9_0 (
            .in0(_gnd_net_),
            .in1(N__2289),
            .in2(_gnd_net_),
            .in3(N__2569),
            .lcout(),
            .ltout(N_90_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIM55C1_6_LC_1_9_1.C_ON=1'b0;
    defparam B_ibuf_RNIM55C1_6_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIM55C1_6_LC_1_9_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 B_ibuf_RNIM55C1_6_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1234),
            .in3(N__2026),
            .lcout(B_ibuf_RNIM55C1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_1_LC_1_9_2.C_ON=1'b0;
    defparam alu_out_RNO_3_1_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_1_LC_1_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 alu_out_RNO_3_1_LC_1_9_2 (
            .in0(N__1974),
            .in1(N__1666),
            .in2(_gnd_net_),
            .in3(N__2290),
            .lcout(alu_out_RNO_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_5_LC_1_9_3.C_ON=1'b0;
    defparam alu_out_RNO_5_LC_1_9_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_5_LC_1_9_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 alu_out_RNO_5_LC_1_9_3 (
            .in0(N__1751),
            .in1(N__1816),
            .in2(_gnd_net_),
            .in3(N__1462),
            .lcout(alu_out_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNII9BS_3_LC_1_9_4.C_ON=1'b0;
    defparam B_ibuf_RNII9BS_3_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNII9BS_3_LC_1_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 B_ibuf_RNII9BS_3_LC_1_9_4 (
            .in0(_gnd_net_),
            .in1(N__2676),
            .in2(_gnd_net_),
            .in3(N__2288),
            .lcout(),
            .ltout(N_87_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIJ25C1_3_LC_1_9_5.C_ON=1'b0;
    defparam B_ibuf_RNIJ25C1_3_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIJ25C1_3_LC_1_9_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 B_ibuf_RNIJ25C1_3_LC_1_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1369),
            .in3(N__2025),
            .lcout(B_ibuf_RNIJ25C1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_3_LC_1_9_6.C_ON=1'b0;
    defparam alu_out_RNO_3_3_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_3_LC_1_9_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 alu_out_RNO_3_3_LC_1_9_6 (
            .in0(N__1504),
            .in1(N__2291),
            .in2(_gnd_net_),
            .in3(N__1667),
            .lcout(alu_out_RNO_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_4_LC_1_10_0.C_ON=1'b0;
    defparam alu_out_RNO_4_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_4_LC_1_10_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 alu_out_RNO_4_LC_1_10_0 (
            .in0(N__1749),
            .in1(N__1837),
            .in2(_gnd_net_),
            .in3(N__1513),
            .lcout(alu_out_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNI6EQF1_4_LC_1_10_1.C_ON=1'b0;
    defparam B_ibuf_RNI6EQF1_4_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNI6EQF1_4_LC_1_10_1.LUT_INIT=16'b0111111100100000;
    LogicCell40 B_ibuf_RNI6EQF1_4_LC_1_10_1 (
            .in0(N__2431),
            .in1(N__1545),
            .in2(N__2307),
            .in3(N__1503),
            .lcout(B_ibuf_RNI6EQF1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIJABS_4_LC_1_10_2.C_ON=1'b0;
    defparam B_ibuf_RNIJABS_4_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIJABS_4_LC_1_10_2.LUT_INIT=16'b0101010110101010;
    LogicCell40 B_ibuf_RNIJABS_4_LC_1_10_2 (
            .in0(N__1546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2278),
            .lcout(N_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_LC_1_10_3.C_ON=1'b0;
    defparam alu_out_RNO_0_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_LC_1_10_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 alu_out_RNO_0_LC_1_10_3 (
            .in0(N__1558),
            .in1(N__1748),
            .in2(_gnd_net_),
            .in3(N__1417),
            .lcout(alu_out_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNI1HJV_0_LC_1_10_4.C_ON=1'b0;
    defparam s_ibuf_RNI1HJV_0_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNI1HJV_0_LC_1_10_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 s_ibuf_RNI1HJV_0_LC_1_10_4 (
            .in0(N__2019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2279),
            .lcout(s_ibuf_RNI1HJVZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_6_LC_1_10_5.C_ON=1'b0;
    defparam alu_out_RNO_6_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_6_LC_1_10_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 alu_out_RNO_6_LC_1_10_5 (
            .in0(N__1798),
            .in1(N__1750),
            .in2(_gnd_net_),
            .in3(N__2686),
            .lcout(alu_out_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam s_ibuf_RNI1PPF_1_LC_1_10_6.C_ON=1'b0;
    defparam s_ibuf_RNI1PPF_1_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam s_ibuf_RNI1PPF_1_LC_1_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 s_ibuf_RNI1PPF_1_LC_1_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2432),
            .lcout(s_c_i_1),
            .ltout(s_c_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIK35C1_4_LC_1_10_7.C_ON=1'b0;
    defparam B_ibuf_RNIK35C1_4_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIK35C1_4_LC_1_10_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 B_ibuf_RNIK35C1_4_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1453),
            .in3(N__1450),
            .lcout(B_ibuf_RNIK35C1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNI08QF1_1_LC_1_11_0.C_ON=1'b0;
    defparam B_ibuf_RNI08QF1_1_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNI08QF1_1_LC_1_11_0.LUT_INIT=16'b0010101011101010;
    LogicCell40 B_ibuf_RNI08QF1_1_LC_1_11_0 (
            .in0(N__1641),
            .in1(N__2478),
            .in2(N__2308),
            .in3(N__1404),
            .lcout(B_ibuf_RNI08QF1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIU5QF1_0_LC_1_11_1.C_ON=1'b0;
    defparam B_ibuf_RNIU5QF1_0_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIU5QF1_0_LC_1_11_1.LUT_INIT=16'b0111111100001000;
    LogicCell40 B_ibuf_RNIU5QF1_0_LC_1_11_1 (
            .in0(N__2479),
            .in1(N__2285),
            .in2(N__1440),
            .in3(N__1960),
            .lcout(un1_A_1),
            .ltout(un1_A_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIE5VR2_0_LC_1_11_2.C_ON=1'b0;
    defparam B_ibuf_RNIE5VR2_0_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIE5VR2_0_LC_1_11_2.LUT_INIT=16'b0111011110111011;
    LogicCell40 B_ibuf_RNIE5VR2_0_LC_1_11_2 (
            .in0(N__2283),
            .in1(N__2020),
            .in2(N__1444),
            .in3(N__1433),
            .lcout(B_ibuf_RNIE5VR2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_0_LC_1_11_3.C_ON=1'b0;
    defparam alu_out_RNO_2_0_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_0_LC_1_11_3.LUT_INIT=16'b0011111001101000;
    LogicCell40 alu_out_RNO_2_0_LC_1_11_3 (
            .in0(N__2480),
            .in1(N__2286),
            .in2(N__1441),
            .in3(N__1961),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_0_LC_1_11_4.C_ON=1'b0;
    defparam alu_out_RNO_0_0_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_0_LC_1_11_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 alu_out_RNO_0_0_LC_1_11_4 (
            .in0(_gnd_net_),
            .in1(N__2201),
            .in2(N__1420),
            .in3(N__1411),
            .lcout(N_142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_0_LC_1_11_5.C_ON=1'b0;
    defparam alu_out_RNO_3_0_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_0_LC_1_11_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 alu_out_RNO_3_0_LC_1_11_5 (
            .in0(N__2513),
            .in1(N__1642),
            .in2(N__2038),
            .in3(N__2287),
            .lcout(alu_out_RNO_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIG7BS_1_LC_1_11_6.C_ON=1'b0;
    defparam B_ibuf_RNIG7BS_1_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIG7BS_1_LC_1_11_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 B_ibuf_RNIG7BS_1_LC_1_11_6 (
            .in0(N__2284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1405),
            .lcout(),
            .ltout(N_85_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIH05C1_1_LC_1_11_7.C_ON=1'b0;
    defparam B_ibuf_RNIH05C1_1_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIH05C1_1_LC_1_11_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 B_ibuf_RNIH05C1_1_LC_1_11_7 (
            .in0(N__2021),
            .in1(_gnd_net_),
            .in2(N__1549),
            .in3(_gnd_net_),
            .lcout(B_ibuf_RNIH05C1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_4_LC_1_12_1.C_ON=1'b0;
    defparam alu_out_RNO_3_4_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_4_LC_1_12_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 alu_out_RNO_3_4_LC_1_12_1 (
            .in0(N__2633),
            .in1(N__2374),
            .in2(_gnd_net_),
            .in3(N__1934),
            .lcout(alu_out_RNO_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_4_LC_1_12_2.C_ON=1'b0;
    defparam alu_out_RNO_2_4_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_4_LC_1_12_2.LUT_INIT=16'b0101111001101000;
    LogicCell40 alu_out_RNO_2_4_LC_1_12_2 (
            .in0(N__2372),
            .in1(N__2482),
            .in2(N__1539),
            .in3(N__1495),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_4_LC_1_12_3.C_ON=1'b0;
    defparam alu_out_RNO_0_4_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_4_LC_1_12_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 alu_out_RNO_0_4_LC_1_12_3 (
            .in0(N__1522),
            .in1(_gnd_net_),
            .in2(N__1516),
            .in3(N__2202),
            .lcout(N_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_5_LC_1_12_4.C_ON=1'b0;
    defparam alu_out_RNO_3_5_LC_1_12_4.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_5_LC_1_12_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 alu_out_RNO_3_5_LC_1_12_4 (
            .in0(N__2375),
            .in1(N__2580),
            .in2(_gnd_net_),
            .in3(N__1496),
            .lcout(alu_out_RNO_3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNI8GQF1_5_LC_1_12_5.C_ON=1'b0;
    defparam B_ibuf_RNI8GQF1_5_LC_1_12_5.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNI8GQF1_5_LC_1_12_5.LUT_INIT=16'b0111001011110000;
    LogicCell40 B_ibuf_RNI8GQF1_5_LC_1_12_5 (
            .in0(N__2481),
            .in1(N__2063),
            .in2(N__1938),
            .in3(N__2371),
            .lcout(B_ibuf_RNI8GQF1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_5_LC_1_12_6.C_ON=1'b0;
    defparam alu_out_RNO_2_5_LC_1_12_6.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_5_LC_1_12_6.LUT_INIT=16'b0101111001101000;
    LogicCell40 alu_out_RNO_2_5_LC_1_12_6 (
            .in0(N__2373),
            .in1(N__2483),
            .in2(N__2070),
            .in3(N__1933),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_5_LC_1_12_7.C_ON=1'b0;
    defparam alu_out_RNO_0_5_LC_1_12_7.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_5_LC_1_12_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 alu_out_RNO_0_5_LC_1_12_7 (
            .in0(_gnd_net_),
            .in1(N__2203),
            .in2(N__1471),
            .in3(N__1468),
            .lcout(N_147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_3_LC_2_9_0.C_ON=1'b0;
    defparam alu_out_RNO_2_3_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_3_LC_2_9_0.LUT_INIT=16'b0011111001101000;
    LogicCell40 alu_out_RNO_2_3_LC_2_9_0 (
            .in0(N__2440),
            .in1(N__2363),
            .in2(N__2677),
            .in3(N__2643),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_3_LC_2_9_1.C_ON=1'b0;
    defparam alu_out_RNO_0_3_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_3_LC_2_9_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 alu_out_RNO_0_3_LC_2_9_1 (
            .in0(N__2198),
            .in1(_gnd_net_),
            .in2(N__1696),
            .in3(N__1693),
            .lcout(),
            .ltout(N_145_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_LC_2_9_2.C_ON=1'b0;
    defparam alu_out_RNO_3_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_LC_2_9_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 alu_out_RNO_3_LC_2_9_2 (
            .in0(N__1861),
            .in1(_gnd_net_),
            .in2(N__1687),
            .in3(N__1782),
            .lcout(alu_out_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNI2AQF1_2_LC_2_9_3.C_ON=1'b0;
    defparam B_ibuf_RNI2AQF1_2_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNI2AQF1_2_LC_2_9_3.LUT_INIT=16'b0111111100001000;
    LogicCell40 B_ibuf_RNI2AQF1_2_LC_2_9_3 (
            .in0(N__2361),
            .in1(N__2438),
            .in2(N__2107),
            .in3(N__1668),
            .lcout(B_ibuf_RNI2AQF1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_2_LC_2_9_4.C_ON=1'b0;
    defparam alu_out_RNO_2_2_LC_2_9_4.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_2_LC_2_9_4.LUT_INIT=16'b0011011011101000;
    LogicCell40 alu_out_RNO_2_2_LC_2_9_4 (
            .in0(N__2439),
            .in1(N__2362),
            .in2(N__1672),
            .in3(N__2106),
            .lcout(alu_out_RNO_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_2_LC_2_9_5.C_ON=1'b0;
    defparam alu_out_RNO_3_2_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_2_LC_2_9_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 alu_out_RNO_3_2_LC_2_9_5 (
            .in0(N__2364),
            .in1(_gnd_net_),
            .in2(N__2647),
            .in3(N__1640),
            .lcout(),
            .ltout(alu_out_RNO_3Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_2_LC_2_9_6.C_ON=1'b0;
    defparam alu_out_RNO_0_2_LC_2_9_6.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_2_LC_2_9_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 alu_out_RNO_0_2_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(N__2197),
            .in2(N__1612),
            .in3(N__1609),
            .lcout(),
            .ltout(N_144_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_LC_2_9_7.C_ON=1'b0;
    defparam alu_out_RNO_2_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_LC_2_9_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 alu_out_RNO_2_LC_2_9_7 (
            .in0(N__1781),
            .in1(_gnd_net_),
            .in2(N__1603),
            .in3(N__1876),
            .lcout(alu_out_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_A_1_cry_0_c_THRU_CRY_0_LC_2_10_0.C_ON=1'b1;
    defparam un1_A_1_cry_0_c_THRU_CRY_0_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam un1_A_1_cry_0_c_THRU_CRY_0_LC_2_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_A_1_cry_0_c_THRU_CRY_0_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(N__1584),
            .in2(N__1588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(un1_A_1_cry_0_c_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_0_LC_2_10_1.C_ON=1'b1;
    defparam alu_out_RNO_1_0_LC_2_10_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_0_LC_2_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_0_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(N__1573),
            .in2(N__1567),
            .in3(N__1552),
            .lcout(alu_out_RNO_1Z0Z_0),
            .ltout(),
            .carryin(un1_A_1_cry_0_c_THRU_CO),
            .carryout(un1_A_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_1_LC_2_10_2.C_ON=1'b1;
    defparam alu_out_RNO_1_1_LC_2_10_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_1_LC_2_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_1_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(N__1912),
            .in2(N__1906),
            .in3(N__1888),
            .lcout(alu_out_RNO_1Z0Z_1),
            .ltout(),
            .carryin(un1_A_1_cry_0),
            .carryout(un1_A_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_2_LC_2_10_3.C_ON=1'b1;
    defparam alu_out_RNO_1_2_LC_2_10_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_2_LC_2_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_2_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(N__2116),
            .in2(N__1885),
            .in3(N__1870),
            .lcout(alu_out_RNO_1Z0Z_2),
            .ltout(),
            .carryin(un1_A_1_cry_1),
            .carryout(un1_A_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_3_LC_2_10_4.C_ON=1'b1;
    defparam alu_out_RNO_1_3_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_3_LC_2_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_3_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__1867),
            .in2(N__2605),
            .in3(N__1855),
            .lcout(alu_out_RNO_1Z0Z_3),
            .ltout(),
            .carryin(un1_A_1_cry_2),
            .carryout(un1_A_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_4_LC_2_10_5.C_ON=1'b1;
    defparam alu_out_RNO_1_4_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_4_LC_2_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_4_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(N__1852),
            .in2(N__1846),
            .in3(N__1831),
            .lcout(alu_out_RNO_1Z0Z_4),
            .ltout(),
            .carryin(un1_A_1_cry_3),
            .carryout(un1_A_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_5_LC_2_10_6.C_ON=1'b1;
    defparam alu_out_RNO_1_5_LC_2_10_6.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_5_LC_2_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_5_LC_2_10_6 (
            .in0(_gnd_net_),
            .in1(N__2047),
            .in2(N__1828),
            .in3(N__1810),
            .lcout(alu_out_RNO_1Z0Z_5),
            .ltout(),
            .carryin(un1_A_1_cry_4),
            .carryout(un1_A_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_6_LC_2_10_7.C_ON=1'b1;
    defparam alu_out_RNO_1_6_LC_2_10_7.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_6_LC_2_10_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 alu_out_RNO_1_6_LC_2_10_7 (
            .in0(_gnd_net_),
            .in1(N__1807),
            .in2(N__2542),
            .in3(N__1792),
            .lcout(alu_out_RNO_1Z0Z_6),
            .ltout(),
            .carryin(un1_A_1_cry_5),
            .carryout(un1_A_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_7_LC_2_11_0.C_ON=1'b0;
    defparam alu_out_RNO_7_LC_2_11_0.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_7_LC_2_11_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 alu_out_RNO_7_LC_2_11_0 (
            .in0(N__2134),
            .in1(N__1702),
            .in2(N__1789),
            .in3(N__1723),
            .lcout(alu_out_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_7_LC_2_11_1.C_ON=1'b0;
    defparam alu_out_RNO_0_7_LC_2_11_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_7_LC_2_11_1.LUT_INIT=16'b0111011110001000;
    LogicCell40 alu_out_RNO_0_7_LC_2_11_1 (
            .in0(N__2122),
            .in1(N__2034),
            .in2(_gnd_net_),
            .in3(N__2128),
            .lcout(un1_A_1_axb_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_7_LC_2_11_2.C_ON=1'b0;
    defparam alu_out_RNO_3_7_LC_2_11_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_7_LC_2_11_2.LUT_INIT=16'b0111000011111000;
    LogicCell40 alu_out_RNO_3_7_LC_2_11_2 (
            .in0(N__2484),
            .in1(N__2379),
            .in2(N__2530),
            .in3(N__2229),
            .lcout(alu_out_RNO_3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_7_LC_2_11_3.C_ON=1'b0;
    defparam alu_out_RNO_2_7_LC_2_11_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_7_LC_2_11_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 alu_out_RNO_2_7_LC_2_11_3 (
            .in0(N__2378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2228),
            .lcout(N_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNII15C1_2_LC_2_11_4.C_ON=1'b0;
    defparam B_ibuf_RNII15C1_2_LC_2_11_4.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNII15C1_2_LC_2_11_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 B_ibuf_RNII15C1_2_LC_2_11_4 (
            .in0(N__2032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2080),
            .lcout(B_ibuf_RNII15C1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIH8BS_2_LC_2_11_5.C_ON=1'b0;
    defparam B_ibuf_RNIH8BS_2_LC_2_11_5.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIH8BS_2_LC_2_11_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 B_ibuf_RNIH8BS_2_LC_2_11_5 (
            .in0(N__2376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2097),
            .lcout(N_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIKBBS_5_LC_2_11_6.C_ON=1'b0;
    defparam B_ibuf_RNIKBBS_5_LC_2_11_6.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIKBBS_5_LC_2_11_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 B_ibuf_RNIKBBS_5_LC_2_11_6 (
            .in0(N__2074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2377),
            .lcout(),
            .ltout(N_89_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIL45C1_5_LC_2_11_7.C_ON=1'b0;
    defparam B_ibuf_RNIL45C1_5_LC_2_11_7.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIL45C1_5_LC_2_11_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 B_ibuf_RNIL45C1_5_LC_2_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2050),
            .in3(N__2033),
            .lcout(B_ibuf_RNIL45C1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_5_7_LC_2_12_0.C_ON=1'b0;
    defparam alu_out_RNO_5_7_LC_2_12_0.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_5_7_LC_2_12_0.LUT_INIT=16'b1110101001000000;
    LogicCell40 alu_out_RNO_5_7_LC_2_12_0 (
            .in0(N__2389),
            .in1(N__2041),
            .in2(N__1978),
            .in3(N__2592),
            .lcout(alu_out_RNO_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_3_6_LC_2_12_1.C_ON=1'b0;
    defparam alu_out_RNO_3_6_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_3_6_LC_2_12_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 alu_out_RNO_3_6_LC_2_12_1 (
            .in0(N__2381),
            .in1(N__2528),
            .in2(_gnd_net_),
            .in3(N__1942),
            .lcout(alu_out_RNO_3Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_2_6_LC_2_12_2.C_ON=1'b0;
    defparam alu_out_RNO_2_6_LC_2_12_2.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_2_6_LC_2_12_2.LUT_INIT=16'b0101111001101000;
    LogicCell40 alu_out_RNO_2_6_LC_2_12_2 (
            .in0(N__2568),
            .in1(N__2487),
            .in2(N__2391),
            .in3(N__2591),
            .lcout(),
            .ltout(alu_out_RNO_2Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_0_6_LC_2_12_3.C_ON=1'b0;
    defparam alu_out_RNO_0_6_LC_2_12_3.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_0_6_LC_2_12_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 alu_out_RNO_0_6_LC_2_12_3 (
            .in0(N__2199),
            .in1(_gnd_net_),
            .in2(N__2695),
            .in3(N__2692),
            .lcout(N_148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNI4CQF1_3_LC_2_12_4.C_ON=1'b0;
    defparam B_ibuf_RNI4CQF1_3_LC_2_12_4.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNI4CQF1_3_LC_2_12_4.LUT_INIT=16'b0111010011110000;
    LogicCell40 B_ibuf_RNI4CQF1_3_LC_2_12_4 (
            .in0(N__2669),
            .in1(N__2485),
            .in2(N__2642),
            .in3(N__2380),
            .lcout(B_ibuf_RNI4CQF1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam B_ibuf_RNIAIQF1_6_LC_2_12_5.C_ON=1'b0;
    defparam B_ibuf_RNIAIQF1_6_LC_2_12_5.SEQ_MODE=4'b0000;
    defparam B_ibuf_RNIAIQF1_6_LC_2_12_5.LUT_INIT=16'b0111000011111000;
    LogicCell40 B_ibuf_RNIAIQF1_6_LC_2_12_5 (
            .in0(N__2486),
            .in1(N__2382),
            .in2(N__2593),
            .in3(N__2567),
            .lcout(B_ibuf_RNIAIQF1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_4_7_LC_2_12_6.C_ON=1'b0;
    defparam alu_out_RNO_4_7_LC_2_12_6.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_4_7_LC_2_12_6.LUT_INIT=16'b0001111011101000;
    LogicCell40 alu_out_RNO_4_7_LC_2_12_6 (
            .in0(N__2529),
            .in1(N__2488),
            .in2(N__2392),
            .in3(N__2230),
            .lcout(),
            .ltout(alu_out_RNO_4Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alu_out_RNO_1_7_LC_2_12_7.C_ON=1'b0;
    defparam alu_out_RNO_1_7_LC_2_12_7.SEQ_MODE=4'b0000;
    defparam alu_out_RNO_1_7_LC_2_12_7.LUT_INIT=16'b1101100011011000;
    LogicCell40 alu_out_RNO_1_7_LC_2_12_7 (
            .in0(N__2200),
            .in1(N__2143),
            .in2(N__2137),
            .in3(_gnd_net_),
            .lcout(N_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // alu_behavioral
